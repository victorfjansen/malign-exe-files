MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ^B*        � �� n   �      }      �    @                      �               @                        �  �	   �   �                   �  �                           �                                                     CODE    Pm      n                    `DATA       �      r              @  �BSS     �   �       t                 �.idata  �	   �   
   t              @  �.tls        �       ~                 �.rdata      �      ~              @  P.reloc  �   �      �              @  P.rsrc    �   �   �   �              @  P             �      6             @  P                                                                                                                                                                �%(�@ ���%$�@ ���% �@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���% �@ ���%��@ ���%8�@ ���%��@ ���%4�@ ���%��@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���%ܠ@ ���%H�@ ���%D�@ ���%@�@ ���%ؠ@ ���%Ԡ@ ��S�ļ�
   T�����D$,t�\$0�Ã�D[Ë��%Р@ ���%̠@ ���%Ƞ@ ���%Ġ@ ���%��@ ���%��@ ���%��@ ���%��@ ��SV�Е@ �> u:hD  j �����ȅ�u3�^[á̕@ ��̕@ 3ҋ���D����B��du���^[Ð� �@Ë�SV���������u3�^[Ë�P�V�P���X�B��^[ËP��
�Q�Е@ ��Е@ �SVWUQ��$��] �$���P�V�;��SS;�u�������C��CF�F;Cu�������CF��;�uË֋��V�����u3��Z]_^[�SVWU����؋��2�C;�rp��J��k;�wb;�u�BC�B)C�{ uH���9����?�΋zϋ�k;�u){�*�
J�$�{{+��|$+��s�ԋ��������u3�����;�u�3�YZ]_^[ÐSVW�ڋ���   }�   �����  ��  ���sjh    Vj ��������;��t#�Ӹԕ@ �l�����uh �  j �P�����3��_^[ÐSVWU�ً���C   jh    h   U�������;��u����  ��  ���sjh    VU������; t#�Ӹԕ@ �������uh �  j �P�b���3��]_^[ÐSVWU���L$�$�D$����3҉T$��$ŉD$�ԕ@ �Q�;�s;�wF��C;D$w;;t$s�t$��C;D$v�D$h �  j V�������u
���@    �������߁�ԕ@ u��D$3҉�|$ t�D$�T$��D$+D$�T$�B��]_^[�SVWU���L$�$�Ћ�� ���$���  �� ����T$�D$�(�D$+ŋT$�B�5ԕ@ �<�^�~�;�v��;|$v�|$;�vjh   +�WS�&�����u
�D$3҉�
�6��ԕ@ u���]_^[Ë�SVWUQ�؋���  �� ����4$���� ����$���+$�A�5ԕ@ �8�^�~�;$s�$;�s��;�vh @  +�WS������u
���@    �6��ԕ@ u�Z]_^[Í@ SVWU��������@ ���?  �� ����] �3;{,�΋׋C�����> tP�FC�F)C�{ u>��������5�;�uɋ֋�������> t!�̋֋�������<$ u��̋V�����3��YZ]_^[Ë�SVWU���$�����@ ���?  �� ����] ��;�t;su�;suW;{��   �L$��+S�CC������|$ t3�L$�T$���]����|$ u��L$�T$�D$�%����$3҉�   �L$�׋������|$ t4�L$�T$�������|$ �f����L$�T$�D$������$3҉�H�k;�u:;{5�$�׋��q����$�8 t(�$�@C�$�@)C�{ u��������$3҉��]_^[ÐSVW�����$���?  �� ����4$��� ���;�s[�ϋ�+Ӌ������L$�׸�@ �]����\$��t�L$�T$���&����D$�D$�D$�D$�|$ t�T$��@ �����3����_^[�U��3�Uh~@ d�2d�"h��@ �9����=5�@  t
h��@ �.����ԕ@ ������@ ������@ �x���h�  j �������@ �=�@  t/�   ��@ 3ɉL��@=  u���@ �@� � �@ ���@ 3�ZYYd�h�@ �=5�@  t
h��@ ������  �堬�@ ]�U��S�=��@  ��   3�Uhb@ d�2d�"�=5�@  t
h��@ �f������@  ��@ P�4���3���@ �ԕ@ �h �  j �CP�%������ԕ@ u�ԕ@ ������@ ������@ �u����̕@ ��t��̕@ P������̕@ ��u�3�ZYYd�hi@ �=5�@  t
h��@ �����h��@ �������!  ��[]�S; �@ u	�P� �@ �P�H��   8;�u��y������@ 3҉T���$��y������@ �T�� ��P[Ë ��P[Í@ ��@ ��J;�rJ;�r����@ u����@    3ҋ�ÐS�ʃ����|�  ����  [Ã�|�ʁ�  ���[����@ �Ѓ�����������@ ��  Ë���|����������Ã�|
�ʁ�  �� ��SV�Ѓ���ʁ�  ���  �t
���@    �ځ����+Ë�3������t
���@    �t �Ѓ��r+�;pt
���@    ����ދ�^[Í@ SVW��3���   �t%����؋�u����X����F�؃#���_^[�SVWU�������$ �������؅���   �k��C�Ѝ7+у���+���+Ń�}�L$��+S׋��������L$�׃��F�����l$��t4��+֋��c�����D$�SS;�s
�7+������T$�������$�$��]_^[Í@ SVW����߉s��ƃ��p��   7�օ�y������@ �D���u��@ �\��[��:��C���Z�,�� <  |�֋��������u� �@ � �@ ��C���Z_^[Í@ �=�@  ~@�=�@ }���@    �+��@ ����@ ���@ ������3���@ 3���@ Ë�SVW������<$���������L$�׸�@ �����\$��u3��R�;�s
����)G�G��t$;�s�����G�G;�u���   ������o���@ �G��@ ���_^[Í@ S����؋ԍC�D����<$ t���W�����u3���YZ[ÐSV�����؋̍V�������<$ t���&�����u3���YZ^[Í@ 3҅�y����=   ��@ �T���u@=  u���SVWU�� �@ ��@ ���@ ;s��   ��C;�~{�s�[;s���B;t��c��   �������؅�uN��������u3��   ;u �)u �} }u 3��E ��@ 5�@ �փ�������@ ��5��@ �L�������S��+ƃ�|��֒�T������;u�C���ƃ ��Ëփ�������@ ��5��@ ]_^[�U����SVW�؀=��@  u	�������t�����~
3��E��T  3�Uh0 @ d�1d�!�=5�@  t
h��@ � ����������}�   ��   ��   �Å�y������@ �T���ty���Ã ��B;�u�Å�y������@ 3��|���&�˅�y�����=�@ �D��
�M��M��A�M���ƋR������E����@ ����@ �  �   ;�@ J)�@ �=�@ }�@ 3���@ ��@ �@ �Ӄ�����E����@ ����@ �A  �2�������E�3�ZYYd�h7 @ �=5�@  t
h��@ �������S  ��E�_^[YY]Í@ U��QSVW��3����@ �=��@  u�f�����u���@    �E�   �a  3�Uh�!@ d�1d�!�=5�@  t
h��@ ����������u���@ 	   ��   ���@ ��%�����)��@ ��tE�ƃ��P��|��  �t���@ 
   �   ��+�;Pt���@ 
   �   ڋ��T����������Ë�;=�@ u,)�@ �@ �=�@  <  ~����3��E���  �   ���t�������}���@    �7��)�ǃx t�8 t�x}���@    ��P�������Ӌ��'������@ �E�3�ZYYd�h�!@ �=5�@  t
h��@ �W�����  ��E�_^[Y]Ë�SVWU�����������}�   ����} �������ǋ�;�u��  ;���   ��+։$;�@ u8�$)�@ �$�@ �=�@ �L  �$�@ �$)�@ ���3  ���u�ËP$������<$|��ދ$����Ã�������   ����   ��+ǉD$;�@ ug��@ ;D$|S�D$)�@ �D$�@ �=�@ }��@ �@ 5�@ 3���@ ��+���@ �E %  ���u ��   �>�������uM�ӋH�$�$;L$}$�ڋ$)D$�,�����D$)$�<$|��Ƌ$�n����:4$��ރ#��.��   �t!%���Ë؋T$���������t	�������3����+���@ �E %  ���u �YZ]_^[Ë�U��QSVW��؀=��@  u�������u
3��E��   3�Uhu$@ d�2d�"�=5�@  t
h��@ �����֋��������t�]��6���������Ã�� %�����;�}�ƅ�t�׋ˑ�b  ��������}�3�ZYYd�h|$@ �=5�@  t
h��@ ������  ��E�_^[Y]Í@ S��~�(�@ �؅�u���   �3ۋ�[�S��t�,�@ �؅�t��   �3ۋ�[Ë��t2��tP���0�@ Y	�t�ð�   ����,�@ 	�u�ð�p   ��tP���(�@ Y	�t�Í@ ��@ �  �SV��؀��=�@  t
�֋���@ ��u��  ��   ���w
3��Ê�4�@ 3��Ë�����^[Ë����$�����PRQ�  ��    YZXu�1������Í@ S���t  ��   [�VW�Ɖ׉�9�wt/��x*�����_^Ít1��|9���x�����������_^�SVWU����S�d����؊��t< v�;"u�{"u����3���C<"u1S�8������S�.�����+��؊��t<"u�; tS�������S������+��؊< w��Ƌ��$  �ߋ>3��Q<"u8S��������S�����;�v��7CF;�w����t<"u�; tS�������S����;�v��7CF;�w��< w���]_^[Ë�SVW�������ڋ����   ��uh  �D$Pj �����ȋԋ���  ��m������Ӌ����������t�; tN���  _^[Ë�SV���f�Cf=��rf=��v�f   �+f=��t���N  f�s�{H u�{ u�CH(@ ���S�؅�t��������^[�f�������Ë�S��3��C3��Cj �CP�CP�CP�P�q�����u�������mu3�[�3�[Í@ 3�ÐSVQ�؋s��u3��&j �D$PV�CP�P�X�����u�����3�3҉SZ^[Ë�S��S�����H��[ÐS��f�C�׋�������u�G���[�3�[ÐV��1��F�Ff�F-��  tHt Ht.�g  �   ��   �   �F�'@ �'�   @�   �   ��   ��   �   �F�'@ �F$((@ �F �'@ �~H ��   j h�   Qj RP�FHP�3�������  �f�~����   f�Nj �6����@��   -�   s1�j j P�6�3���@��   j ��j Rh�   ��L  R�6�����ZH��   1�9�sk��L  t@��jj )�P�6�����@��   �6�����Huv�=��L  �F�   �F$�'@ �Ff�~��tj����Г@ uj��j��x������t9�f�~��t�6�R�����t��u�F �'@ 1�^��6�'���f�F�׸i   ��f�F���������SV��؋�3ɺL  �   ��L  �Cf�C��3���@ f�C�C�   �CH(@ ���-  P���%  �SHY�d������  �DH 3�^[Í@ Sf�Hf���tIf��s���Ӌ��3��=�@ t=Г@ u3���g   ��t���������[Í@ �P ����Í@ SV��3�f�Cf=��r/f=��w)f%��f=��u���S����u���S$����t���������8�@ t
�g   ������^[Ë�W�ǈ͉���f�ȉ���x	�у��_ÐSVW��P��tl1�1ۿ����F�� t�� ��-tb��+t_��$t_��xtZ��XtU��0u�F��xtH��XtC��t ���t-��0��	w%9�w!���؊F��u���t	��}T�	F���~KxI[)��G�ŊF뜿����F��t߀�ar�� ��0��	v����wЀ�
9�w���؊F��u���u��Y1��2_^[Í@ S�؁��@ t��Г@ u3���@ f�C���o���f�{�����؄�u
�i   �b�����[Ë�VW��f�x��tPRQ������YZXt5�xx�P+P9� P)�PQ����P��uYX������YX_^�H�_^Ð�Ѻ�,@ ��@~d��@PQ�@   �����d  ��    uYX��YX�                                                                ���4���Í@ SVQ���Ct�$�D$
�ԋù   ��������$
�ԋù   ����������S�����Z^[Ð�%0�@ ��S3�j �������uj�����% �  =   t=   u���[ÐU������@ �E��E�Pjj h(.@ h  �������uM3�Uh.@ d�0d� �E�   �E�P�E�Pj j hD.@ �E�P�����3�ZYYd�h.@ �E�P������  ��f��@ f%��f�U�f��?f�f��@ ��]� SOFTWARE\Borland\Delphi\RTL FPUMaskValue    ���-�@ Ë���t���Q�À=�@ vj j j h�����@ Ð�=�@  tPPRTjj h�����@ ��XÍ@ Tjj h�����@ ��XÍ@ �=�@ vPS�����Í@ ��t�A�9�t�9�u��AA����Ë��=�@ vPRQ�����QTjj h�����@ YYZXÐ�=�@ vRTjj h�����@ Z�PR�=�@ vTjj h�����@ ZXË��D$�@   �  �8����P�Htn��������@ ����   �҅���   �T$�L$�9���t7������=�@  v)�=�@  w �L$PQ������ X��   �D$�H�0�D$�H�=�@ v�=�@  wP�D$RQP�H����� YZXtp�HS1�VWUd�SPRQ�T$(j Ph40@ R��@ �|$(��  ��    ��    �o�_�G`0@ ���f������#   �  ��    ���    �A������   Ë��D$�T$�@   t�J�B�0@ SVWU�j���F�����]_^[�   Ë��D$0�@1@ �H  ��    �
��    �B�`��8���t�B�k����r���1���d�Y��]_^[�   Í@ ��  ��    �
��    �B�1���Z�d$,1�Yd�X]��������1ҋL$�D$��d���� Ë�U��U�=�  �,t\=�  �tW-  �t\-�   t=HtN�`q��?��r6t0�R=�  �t=-�  �t.HtHt$�:-�  �t/��=t&�,���*���&���"������������������
��������%�   �R� ���]� �D$�@   ��   �=�@  w�D$P�0����� tq�D$��%����T$j PhB2@ R��@ �\$�;����S�Ct��@ ����������҅�������S�������@ ��t�ыL$��   �Q�$�J  1�Í@ 1ҍE�d�
d���@�1@ �h�$�@ Í@ 1ҡ$�@ ��td�
9�u� d�Ë	���t9u�� ��U��SVW� �@ �G��tH�_�p3�Uh*3@ d�2d�"��~K�_�D���t�Ѕ��3�ZYYd���-����������������_^[]ÐU��SVW�(�@ ��tK�03ۋx3�Uh�3@ d�2d�";�~��C�,�@ ��t��;��3�ZYYd��������P����'����v���_^[]Ð��@ (@ ��@ 8@ �(�@ 3��,�@ �0�@ �B��@ ������$�@  �a����SVW�X�@ �� �@ �ÿ
   �����03�����û
   �����I��u۱��@ �Ѓ���x�@ 3ۊو��I��u�_^[Ë�1�� �@ ���@� �@ �_�o�w�w �7�   �_^�� Ë�Q�=4�@  tWf�=�@ ��u�=�@  v��@ � �@ j �D$PjhX�@ j��r���P����j �D$Pjh�4@ j��W���P����ZÀ=�@  uj hP�@ hX�@ j ����Z� ����   
  SVWU� �@ � �@ �0�@ �{( u�? t���3҉���Ճ? u�=�@  t�����2���3���@ �{(u
�> u3��C�����{(v�> t!�C��t�#  �S�B;Bt
��tP������1����{(u�S$�{( t�����; u�=�@  t��@ �P�����V�����   �^�v���]_^[ã �@ ����Ð��@ �����Ë��t�     �J�I|��J�u
P�B�����XÐSV�É֋��t�    �J�I|��J�u�B��r�����Nu�^[Ð��t$�J�APR�B��\   ��XR�H��L���ZX���B����t�J�I|��J�u�B��&���Ð��t
�J�A~��B����t�J�I|��J�u�B������Í@ ��~$P��
���P�����Zf�D�  ��Z�P��@�   �1�ÐSVW�É։ω���������ǅ�t	��������������;_^[Ë�R��   �����ZÐ1Ʌ�t!R:
t:Jt:Jt:Jt����BBB��Z)�����Í@ WPQ��1��u��X�X_�y���Å�t�@�Å�t?��������SVW�É֋y��V��9�t�  ���N�������_^[���  �����Å�ta�������;t\;tPQ�u���ZX����SVW�Ӊ�P�C�F�������ǉ؋K����������N�S�����X����t�O��/���_^[É��$������I����SVWRP��1��L���t9u�ϋA�J�1��L���t	A�9�u1�Ju��t�$�w��,  �<$�77K��9���P�ƋD����t
�H������Ku�ZX��u��t�J�����Z_^[X�$���Ë�SVW�Ɖ�9���   ��th��tk�F��W�)�w�R��t&��9�uXJt�N�_9�uK����Ju������Z��t"��8�uAJt8�u:Jt��  � ��  � 9�u'��#�W�)���F�)��Z8�u8�u����8�u8�_^[Ë���t
�P�B~��@�Ð��t� �i9@ Ë��t8�J�It2S�ËB��)�����P�H�����X�H�I|��H�u�@�������[��Í@ ����Ë�����Ë�S��t-�X���t&J|9�})Ӆ�|9�D$������1������D$�����[� �SVW�É։��������t0�J�N|*9�}&��~")�9�~��)���r�����؋R�)��L   _^[Å�t@��t1SVW�Ɖ׋O�W�V�Jx�F)�~�u��VW���_^t����Z1��1��Z��)�_^[Í@ SVW�É�1���~H���t#�x�u����	P������X����p�� �(��������ǋ��t���H�9�|���������������;_^[Ë�3��   �S�Ӊ�1Ʌ�t�K�)�Q�~���Y��[�!���ð�I����U����SVW�E��$�@ �E��}� t93�Uhc;@ d�0d� �]��E��S3�ZYYd��
����������E�� �E��}� u�_^[YY]Ë�� �@ �� �@ Ë�U��Q�E�3�Uh�;@ d�2d�"�E��@�t���3�ZYYd�h�;@ �E�; �@ u�E�� � �@ �� �@ ��t�;U�u	�U����� ��u��������Y]Ë�U����S3҉U�3�Uhj<@ d�2d�"j�U�Rh  P�a����E��U��   �����E��U�������؃}� t3�3�ZYYd�hq<@ �E��������������[��]�U��3�Uh�<@ d�0d� ���@ u#�8�@ ������@ �����Г@ ���������3�ZYYd�h�<@ ��������]Ð�-��@ ��   ��@ ��@ (@ ��@ 8@ �6�@ � �@  ;@ �V�����t�}����<���f�<�@ ��f��@ ��f�ԓ@ ���H����,�@ �����(�@ ����%   �=   �t-�s���%�   f��v���@    � �/����������@ ������u������@ �/���� �@ Ð�%\�@ ���%X�@ ���%T�@ ���%P�@ ��Pj@�����Í@ �   Ë�S������؅�t6�=��@ �u
��   ��������������u��   ������P���@ P����[ÊL�@ ���@ ��u&d�,   ����������@ P�n�����táX�@ �P�]�����t�ø��@ �"���ÐS��3����@ j �+����P�@ �P�@ ���@ 3����@ 3����@ ��������@ ������[Í@ U��3�Uh�>@ d�0d� �T�@ 3�ZYYd�h�>@ �������]Ë��-T�@ �U��3�Uh?@ d�0d� �\�@ 3�ZYYd�h?@ ��~�����]Ë��-\�@ ��%l�@ ���%h�@ ���%d�@ ���%<�@ ���%8�@ ���%4�@ ���%0�@ ���%,�@ ���%(�@ ���%$�@ ���% �@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���% �@ ���%��@ ���%��@ ���%��@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���%ܡ@ ���%ء@ ���%ԡ@ ���%С@ ���%̡@ ���%ȡ@ ���%ġ@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%|�@ ���%x�@ ���%t�@ ���%`�@ ���%\�@ ���%X�@ ���%T�@ ���%P�@ ���%L�@ ���%H�@ ���%D�@ ��U�����U��E��E�3ɋU������YY]Í@ U�����E�3��E��E�YY]Í@ U��3�UheA@ d�0d� �`�@ 3�ZYYd�hlA@ �������]Ë��-`�@ ��%l�@ ���%h�@ ��U��3�Uh�A@ d�0d� �d�@ 3�ZYYd�h�A@ ��������]Ë��-d�@ �SV��؋�����P������P������P������Pjh   �F�����^[�SVW�������^����؃�|(�D�</t<\t<:uW�S�����������K��}؋ǋ�����_^[Ë�SV��؋Ƌ������^[Ë�SVWU������������   �C;�|�|� v�;�}
���e����N�|7� v�U��+�A�Ӌ��$���]_^[Í@ U��Ĵ���S�؍�����P������P��������t4P�����������u%�E�P������P�����E�P�E�P�E�P������u�E������E�[��]�S�؋�����@��[�SVW�ڋ���������w?�Ӂ��   ��@w2j h�   jj ��%�   ������@ P����@ P�������P�����_^[ÐQj RP�����ÐSVWQ�����j �D$PWVS������u�$�����$Z_^[�P�z���ÐS�؋�����P�������t�u3�[ð[Í@ U��3�UhD@ d�0d� �h�@ 3�ZYYd�hD@ �������]Ë��-h�@ Ã��3ɉ$�L$Q�L$Qj h?  j j j RP������$YZÉ��ǹ����2������)ȉ�ÐU��QSV�M��u�����؋������PVjj �E�PS����S����^[Y]� �U��3�Uh�D@ d�0d� �l�@ 3�ZYYd�h�D@ ��������]Ë��-l�@ �U��QSVW�E��E��z���3�Uh�E@ d�0d� 3�Uh�E@ d�0d� �x�@ ������t!�   �x�@ �����ع   3ҋ��U����
3�ZYYd��_���u
3�ZYYd��P�u�h�E@ h�E@ �E��   ������E�����P�E��S����Ћ�Y�������6���3�ZYYd��
���������3�ZYYd�h�E@ �E��I�����������_^[Y]�   ����      ����   
   U��3�QQQQ3�Uh�F@ d�0d� �U���F@ ��  �U��p�@ �C����U���F@ �  �u��5p�@ �U���F@ �  �u��x�@ �   ������U��F@ �q  �U�|�@ �p�@ �^����t�@ �p�@ ��F@ �I���3�ZYYd�h�F@ �E�   ������������]�   ����   ��  ����   ú����� ����   ����    ����   ��������    ����   r   U��M�A��E�P�]Í@ U��QSVW�M�����3ۋE�PWV�����U�B�E�x� tC�E�@�PV�)����U�B��E�x� t'�EP�E�@�PV�I���P�E�@�P����Z����Y���_^[Y]Í@ U����SVW�M�U�E�E�������E�������E������3�Uh�H@ d�0d� U�E�����P�E������СP�@ Y�1���Y����   �E��@�����t�E�����P����3�UhjH@ d�0d� j h�   jj j h   ��E��Z���P�@����؀} t.�E�Mj �E�Pj�E�PS����j �E�P�E�HP�E�@PS�t����j �E�P�E�P�E�PS�^���S�����3�ZYYd��
����������E������E�P�3���3�ZYYd�h�H@ �E�   �q�����������_^[��]� U����SVW3ɉM���E��E�����3�Uh:I@ d�0d� �������E��|�������~.�E�   �E��U��\��À�E��� ����U���V����E�Nu�3�ZYYd�hAI@ �E������E�������I�����_^[��]�U����SVW3ɉM�U��E��E������3�Uh�I@ d�0d� �E��r����E����������~B�   �E��\0���%  �yH���@��u��9���&�E���T����U�E������E�FOu�3�ZYYd�h�I@ �E������E������������_^[��]Ë�U��3�UhGJ@ d�0d� ���@ u(�|�@ ������x�@ ������t�@ �����p�@ ����3�ZYYd�hNJ@ ��<�����]�U��SVW3�Uh�J@ d�0d� �-��@ s'3�Uh�J@ d�0d� �L���3�ZYYd��
���������3�ZYYd�h�J@ ��������_^[]Ë�U��3�QQQQQQQS3�Uh1L@ d�0d� �=��@  �&  h@L@ �������@ �=��@  �
  �U��XL@ �����E��[���P���@ P��������@ �U��|L@ �����E��5���P���@ P�������@ �U���L@ �c����E�����P���@ P�������@ �U�L@ �=����E������P���@ P�i������@ �U��L@ �����E������P���@ P�C������@ �U��L@ ������E�����P���@ P�������@ �U��L@ ������E��w���P���@ P��������@ �=��@  t	�=��@  u3���3�ZYYd�h8L@ �E�   �������R������[��]� kernel32.dll    ����   ����������������������    ����   ������������  ����   �����������   ����   �����峲�����   ����   �����峲����    ����   �����䳲�����   ����   �����䳲����    SV���������tVS���@ ^[�3�^[ÐSV���������tVS���@ ^[�3�^[ÐSV����a�����tVS���@ ^[�3�^[ÐU���D�����t�EP�EP���@ �3�]� ��U��� �����t�EP�EP���@ �3�]� ��U��3�Uh�M@ d�0d� ���@ 3�ZYYd�h�M@ �������]Ë��-��@ �U��hN@ hN@ �2  �P���UR��]� GetCurrentThreadId  Kernel32.dll    U���d���SVW�}�]ǅd����   ��d���P�����j2�%�����t���uWS��   �   �[���P�i����E�S�`�����j`S������t3��   �;t3��   �C8P�6���������;�u	�
������Vj h� ��������u3��Tj Wh� �E�P�����PjV�����������;�tV�,������@��u3���E����U��RD��Ѓ���E�_^[��]� ��U��j j S3�Uh�O@ d�0d� �U��P@ �U����E�����P�������@ �U��P@ �5����E������P��@ P�a�����@ �E��@ �E�Ԁ@ h��@ hȀ@ h� hĀ@ ��@ ��@ P������Ā@ 3�ZYYd�h�O@ �E��   �'�����������[YY]�   ����	   ��������   ����   ������������    U��S�EP�����؅�u3���EPS�����Ѕ�u3���8huB�[]� SVW����3���3ɺ   ����3Ҹ   �����؃��t/�$   TS�������t;|$u�t$�TS�������u�S�v����ƃ�_^[ÐU��3�Uh�P@ d�0d� ���@ 3�ZYYd�h�P@ �������]Ë��-��@ øj ��3���t��Í@ U��SVW�؅�tB3�UhRQ@ d�2d�"��f�8�%u�@��À8hu	�x�u�X3�ZYYd������3�������_^[]Í@ U����SVW3҉U�U���3�Uh�R@ d�0d� 3۾Q@ ���P@ Wj h� ��������@ �=��@  ��   j@h   Vj ���@ P��������@ �=��@  ��   �U�R@ ������E��s���P������؍U��R@ �����E��V���PS�����������E�Vj �����؅�tT�Ӹ�P@ ���s����փ���| B�E�    ��E��8u�M��E�Ju�E�PVS���@ P���@ P�G���S�����3�ZYYd�h�R@ �E�   �u������������_^[��]�����   �����쳲����    ����   ����������� SVW��4�����3�j V�?������@ �=��@  tu�=��@  tl���@ P�����$  T���@ P�������t1V�t$���@ �3   �^���@ ��$�   �$  T���@ P�1������@ P����j j j V������Á��   _^[�SQ���$ ��t'���������t��������؅�t���1�����t�$�$Z[Í@ U��3�Uh�S@ d�0d� ���@ 3�ZYYd�h�S@ �������]Ë��-��@ �U��   j j Iu�Q3�Uh�T@ d�0d� �U��U@ �����E��A���P�U�� U@ �����E��+���P����j j jP�����U��4U@ �X����E��  �U�U@ �C����E��  �U�HU@ �.����E��n  �U�\U@ �����E��Y  �U�pU@ �����E��D  �UคU@ ������E��/  �Uܸ�U@ ������E��  3�ZYYd�h U@ �Eܺ	   ������������]�����
   ���������  ����   ����������� ����   ���������� ����   ������Ү��� ����   �������    ����
   �����Ԯ���  ����   ������ή��� ����
   �����׮���  U�������SVW3҉������������������E��E�����������3�Uh�V@ d�0d� 3�3Ҹ   �������(  �׋��"������@�n�������W$�  �/���������������������������U�������t%�������W$�  ������������U��_�����u���׋���������@��u�V����3�ZYYd�h�V@ �������   �q����E��E�������������_^[��]�U����SVW3ɉMȉM̉U��E�3�Uh�W@ d�0d� 3��E�U̸�W@ ������E��m���P�K����؅�tr�Uȸ�W@ �����E��L���PS�����������tN�E��E�3��E��E�   3��E�3��E�3��E�3��E�3��E�E�P�E�P�E�P�E�P�օ�t3��E���E��E�3�ZYYd�h�W@ �EȺ   ������������E�_^[��]�   ����	   ��������   ����   �������������   ��l����$�   T�=����|$u3����Ĕ   ÐU�������SVW3҉������������������������E��E��+���3�Uh�Y@ d�0d� 3���3Ҹ   ������ǅ����(  ����������������@�,  �������������  ������������������f����������U�� �����t,�������������  �����������U����������   ������Pj�j�����؅�tL��u.��������Y@ �����������_���Ph�Y@ �8���P���������tj S�׃��@�E�S� �����E� �}� uH������u?�������   �c����؅�t)��tj S�׃��@�E�S�����}� u��������������������������@�������V����3�ZYYd�h�Y@ �������   �N����E��"����������_^[��]�   ����   ����������������    kernel32.dll    U��3�Uh-Z@ d�0d� ���@ 3�ZYYd�h4Z@ ��V�����]Ë��-��@ Á�l����$�   T������|$u3����Ĕ   ÐSV��  �Ƌ�����S���:���P�����؋Ƌ�������|�\t�ƺ�Z@ �����^[� ����   \   SV��  �Ƌ������S�������P�(����؋Ƌ�������|�\t�ƺ[@ �t���^[� ����   \   U��3�Uh-[@ d�0d� ���@ 3�ZYYd�h4[@ ��V�����]Ë��-��@ �U��İ���S3��������������������������������������������������������E�3�Uh�]@ d�0d� ƅ���� ������Ph  �e���ƅ���� ������Pj h�]@ ������P�<�����������]@ �����������P�������������P����������E�Y�����E��Y�����S�]����U���(����������(����d����K�����������]@ �o�����������(������������ ���h ^@ ������3��j���������h^@ �������   ������������(����^����q��������h^@ ������3��"���������h^@ �������0^@ ������������������   �=�����������(���� ��������z���h ^@ �u�h^@ �������   ������������(��������������B�����(����k����2���������3ɺD   ����ǅ����D   ǅ ���   fǅ���  �����P������Pj j j j�j j Sj �������3�ZYYd�h�]@ �������	   �V����E��*�����������[��]� $$cd    ����   ����    ����   ����    ����   del "   ����   "   ����
   if exist "  ����	   ��������   U����S3҉U��E��E�����3�Uh�^@ d�0d� 3ۍU���^@ �@����E��U�������E������Pjj j ��������@ �=��@  t�>���=�   u�3�ZYYd�h�^@ �E��   �K�����������[YY]�����   �����   U��*   j j Iu�SVW��3�Uh.b@ d�0d� �������Db@ ������������������  �E�Pj �D�����u�E�j j �;�����E� k�����  @�E��E��Tb@ ����j hdb@ �u�hpb@ �������   �������������������������������P�(���������  3۾   �E���b@ ����j hdb@ �u�h�b@ �������   �?��������������������������c���PSW������؅��  h   ������PS����Ƅ���� �������������   �	���������P��������b@ �V���������X�J�����   �������������   �����������P��������b@ ����������X����t}�������������   ����������P��������b@ �����������X�����tB�������������   �T���������P��������b@ ����������X����tN�������tj j h�   S������H3۾   j ��������b@ �^�������������PSW�s����؅�tNu҅�tj j h�   S�w����E���b@ �����j hc@ �u�hc@ �������   �w������������������������������P��������tj j jW����jd�����M��i����}� t�}� t�E�Pj �x���3�ZYYd�h5b@ �������   ������E�������U�����_^[��]�����   ������ ����   Ю��    ����   ��  ����	   ���������   ����   Ю��    ����   ����    ����   TJPm    ����   Lx9}    ����   $93�    ����   8u9�    ����
   ��Ю������  ����   ��������    ����   ��Ю    ����   ������������    U��
   ����3�]� �U��ĨS�ډE��E�� ���3�Uh�c@ d�0d� �E��D   �����E�D   ��u�]�S�E�Pj j j j�j j �E������Pj ��������@��3�ZYYd�h�c@ �E��1�������������[��]Ë�U��QSVW�E��E��v���3�Uh8d@ d�0d� 3��E��n����؅�y����K��|C3��E���������B�D�8FKu�3�ZYYd�h?d@ �E�������K�������_^[Y]ÐU��   j j Iu�3�Uh�e@ d�0d� �E���e@ �����E���e@ �U��.����E�U��#����U����@ �����E���e@ �����h�e@ �u�h�e@ �E�   �c����E�U�������U𸘗@ �g����E���e@ ����h f@ �u�hf@ �E�   �$����E�U������U踠�@ �(����E��f@ �_����Eܹ8f@ �U��{����E܍U��p����Uฐ�@ ������Uظ\f@ �V����M؋�@ ����@ �A���3�ZYYd�h�e@ �Eغ
   �������������]�   ����   ����    ����   ��������    ����   ����    ����   ��  ����   ������  ����   ����    ����   ��  ����   ������  ����   ������������������  ����   ��������������������������� ����   ������  U��Q�H   j j Iu�Q�M�SVW�M�U��E��E�������E�������E�����3�Uh
i@ d�0d� ��E�M�U�������E�M�U�������E��@�����u3��  �E��-�����uj �E��s���P�E��j���P�@����E������h�  ����j �E��H�����V������3�謿���������-���P��������  �E�$i@ �U��[���j �E�����P������3��k��������������P��������Y  �E�x� ��   h  ������P�E�����P�K���h  ������PV�9����������4i@ ���������������P�h������������Li@ �����������g���PW��������������pi@ �����������C���P������P������P��������i@ �p�������������P���   �E�����h�  �3���j V������3��c��������������P������uU�������4i@ ��������������P��������������i@ ���������������PW�!�����jV�E�����P��3�ZYYd�hi@ �������	   �����E�   ������y����ۋ�_^[��]�  ����   .ddd    ����   �����̳�����    ����   ��������������������������  ����   ����������� ����   ������  ����   ����������� U��   j j Iu�SVW3�Uho@ d�0d� �Uܸ0o@ ������E������E�������E�P�   �   �E�������E�P�UԸ<o@ �����MԍE�Z�����U�3�込���EЍU���������@ �E�������t(���@ �E��{�����t���@ �E��i�����t3���������E��}� tO�U̸To@ �4����E������P�������Uȸlo@ �����E������PV�H�������t
j����P��V������]��  ������ЍE��F����EčU��w����E�P�   �   �E�������E���o@ ����u1�E��   �   ������U���o@ �'����H�E��   ������+�U���o@ ������u
�E�������U��ȸ   ��������@ �E��P�����u/h�o@ �u��5��@ h�o@ �u��E��   �����E�3������?���@ �E�������u-h�o@ �u��5��@ h�o@ �u��E��   �L����E�3��^�������  �}� tF�}� tU���@ �U܋E��\���Y�U���@ �U܋E��G���YU���@ �U܋E��4���Y�H  �E���o@ �A���h�o@ �u�h�o@ �E��   ������E��U��H����E������E���o@ ����h�o@ �u�h�o@ �E��   �����E��U������E��N����U��p@ ������E��9����U��p@ ������M��E��U�������E��������uj �E��t���P�R����E���@ �U�����j �E��S���P�U�3�輹���E��@���P��������   ���@ ǀ]     ����@ P�����h�  �@������@ �������uݡ��@ P����j j jh��  �w���h�  �������@ 3҉�]  j �E������P�U�3��+����E�����P�����U��,p@ ������E�����P�U��To@ ������E��~���P�\���P������ÍE�Pj j h,c@ j j ��h�  �����E��K���P��@ � �>���P���@ �3����и  �Y�����= �@  t7���@ P��������@ P�K������@ P����������3ҋE������j �������@ ������tf���@ P�������@ ǀ]     ����@ P�}���h�  ��������@ �u�����u�j j jh��  ����h�  �������@ 3҉�]  3�ZYYd�h!o@ �E��   �����E��   �������i�����_^[��]�����   �� ����   �������������  ����   �����̳�����    ����   ����������������������  ����   "   ����       ����   "   ����   ��  ����   ����    ����   Ю���   ����   ����    ����   ��  ����   ����    ����   ���Ю���    ����   ������  ����   ������������    U��   j j Iu�SVW���@ 3�Uh�s@ d�0d� ��@ � �����Ph.]  j jj j���������@ j j j j���@ P��������    �3҉�]  �3҉�!]  �3҉�]  ����@ ��)]  ��@ ���-]  ǅ@����   ��@���P�/�������������E�s@ �|����E�������t
�H���������3҉�]  ��<����@x@ �x�����<�����@ ��E��b�����8����_�����8����E�M��F����E�������t�E������P�����j��4����Px@ ������4���P��0����`x@ ������0����M�Z�����E�����P�~����؅�u�E�����P�j����؅��s  ��,����lx@ ������,����a���PS������Ǎ�(����xx@ ������(����=���PS������E��� ����|x@ ������ �����$����^�����$��������؋E�������Ѝ�����������������������������E���������@ P�����P�   �   �E������������{@ �������PS�����P�����   �E������������y���P�׋3҉�]  ���]  tFjj j j �E�P�������t�}�t+�E�P������E�P����h�  �^����������!]  ��U�h   h��@ ����3�ZYYd�h�s@ ������   �����E�   ������������_^[��]������  JiF����sUh������T������g���h��U����g���x������c���fj\lT���L��������v ***/2;********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************* 	 ����   ������ ����   ���    ����   ��� ����   �  ����   �   ****************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************  ����   $   U��3�Uh�{@ d�0d� ���@ u2���@ �E������@ �;������@ �1������@ �'������@ ����3�ZYYd�h�{@ �馴����]Ë�U��3�Uh)|@ d�0d� �-��@ s�<|@ �����7����<|@ ����3�ZYYd�h0|@ ��Z�����]�  ����'                                           U��3�Uh�|@ d�0d� 3�ZYYd�h�|@ �� �����]�   �|@ �>@ �>@ �<@ x<@ ?@ �>@ pA@ @A@ �D@ �D@ D@ �C@ PJ@ �I@ �M@ �M@ 8[@ [@ �P@ �P@ �S@ �S@ 8Z@ Z@ �A@ �A@ �{@ �{@     d|@ U����SVW��|@ �E���3�Uh<}@ d�0d� �
���3�ZYYd��
�����γ��_^[讷����                                                                                                                                                                                        �@ 2�� �@  �@  �@ �@         �@ D @ �#@  ��������������������� ��@ Error ��Runtime error     at 00000000 ��0123456789ABCDEF����                           �   @   �                                                               ��VqDR3          |�@ p�@ t�@                                                                                                                                                                                                                                                         t�  ��              ��  0�              ��  @�               �  P�              L�  d�              ��  t�              �  D�              ��  h�                      ��  ��  ��  ʢ  �  ��  �  �  �  ,�  B�  T�  f�  |�  ��  ��  ��  ��  ̣  أ  ��  �  �  "�  .�  @�  P�  ^�  l�  z�      ��  ��  ��      Τ  �  �      �  �  *�  8�      Z�  l�  ~�      ��  ��  ��  Υ  �  �  ��  
�  �  .�  @�  P�  ^�  n�  ~�  ��  ��  ��  ��  ʦ  �  �  �  �  *�  @�  T�  f�  z�  ��  ��  ��  ʧ  ܧ  �  ��  
�  �  (�  B�  Z�  h�  z�  ��  ��  ��  Ĩ  Ҩ  �  �  �      �  2�  B�  X�  h�  z�  ��  ��      ��  ʩ      kernel32.dll    DeleteCriticalSection   LeaveCriticalSection    EnterCriticalSection    InitializeCriticalSection   VirtualFree   VirtualAlloc    LocalFree   LocalAlloc    GetVersion    GetCurrentThreadId    GetThreadLocale   GetStartupInfoA   GetModuleFileNameA    GetLocaleInfoA    GetLastError    GetCommandLineA   FreeLibrary   ExitProcess   WriteFile   UnhandledExceptionFilter    SetFilePointer    SetEndOfFile    RtlUnwind   ReadFile    RaiseException    GetStdHandle    GetFileSize   GetFileType   CreateFileA   CloseHandle user32.dll    GetKeyboardType   MessageBoxA   CharNextA advapi32.dll    RegQueryValueExA    RegOpenKeyExA   RegCloseKey kernel32.dll    TlsSetValue   TlsGetValue   LocalAlloc    GetModuleHandleA  advapi32.dll    RegSetValueExA    RegCreateKeyExA   RegCloseKey kernel32.dll    WriteProcessMemory    WriteFile   VirtualAllocEx    UnmapViewOfFile   SuspendThread   Sleep   SizeofResource    SetThreadContext    SetLastError    SetFilePointer    ResumeThread    OpenProcess   MapViewOfFile   LockResource    LoadResource    LoadLibraryA    IsBadReadPtr    GlobalFree    GlobalAlloc   GetWindowsDirectoryA    GetVersionExA   GetThreadContext    GetTempPathA    GetTempFileNameA    GetSystemDirectoryA   GetShortPathNameA   GetProcAddress    GetModuleHandleA    GetLastError    GetFileAttributesA    GetCurrentProcessId   GetCurrentProcess   GetCommandLineA   FreeResource    FreeLibrary   FindResourceA   FindFirstFileA    FindClose   FileTimeToLocalFileTime   FileTimeToDosDateTime   ExitProcess   DuplicateHandle   DeleteFileA   CreateSemaphoreA    CreateProcessA    CreateFileMappingA    CreateFileA   CreateDirectoryA    CopyFileA   CompareStringA    CloseHandle user32.dll    TranslateMessage    SendMessageA    PostThreadMessageA    PeekMessageA    GetWindowTextA    FindWindowExA   FindWindowA   DispatchMessageA  winmm.dll   waveOutSetVolume    waveOutGetVolume                                     �@ �@ ��@ �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ,  0
000"0*020:0B0J0R0Z0b0j0r0z0�0�0�0�0�0�0�0�0�0�0�0�01111&1.161?1`1h1�1�13�3�3+4>4�4�495m5y5�5'6v7�7�7�7�7�7�788!8'858H8R8X8f8l8t8�8�8�8�8�8�8�8�8�8�8�8999$9/9@9F9N9X9o9z9�9�9�9�9�92:H:�:�:�:�;<?<E<^<g<p<{<�<�<�<�<�<=$=�=�=�=�=>>D>T>]>�>�>�>�>�>�>.?X?r?�?�?�?�?�?�?�?�?�?�?�?      �   00&0P0V0h0�0�0�0�0�0�0�01&1.141:1l1�1�1�1�1�112<2E2K2[2d2�2�2�2�2�2�2�2�2�23�3�3�3�34]4c4k4�4�4�4�4	55/5<5\5u7{8�8�8�8�9�9�9:,:|:�:�:<	<<�<Z=�=�=�=�=�=
>>Y>n>�>�>�>�>�>�>?"?6?@?S?�?�?�?�?�? 0  (  )000R0�0�0272>2V2x2�2�2�2�2 3K3^3r3�3�3�3�3�3�3�3�3�3�3�34'4D4N4s4}4�4�4�4�4�4�4�4�4555-5A5�5�5�5�5k95;F;�;�;�;�;�;�;�;<]<<�<�<�<�<�<�<�<�<�<�<�<�<�<==$=-=9=C=j==�=�=�=�=�=�=�=>>>8>H>Y>j>v>{>�>�>�>�>�>�>�>�>�>�> ???"?*?2?:?B?J?R?Z?b?j?r?z?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   @  0  0
000"0*020:0B0J0R0Z0b0j0r0z0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01G1S1`1r1z1�1�1�1�1�1Y3a3�3�3�34�4�4�4�4�4�4�4
5B5G5�5�5�5�5666$666C6I6S6Y6^6p6�7�7�7�8�8%9h9�9�9:::&:0:B:Z:f:q:�:�:�:�:�:�:�:;;;1;<;D;W;b;j;};�;�;�;�;�;�;�;�;�;�; <	<<=7=W=z=�=�=�=�=�=�=�=D?R?j?r?�?�?�?�?�?�?�?�?�?�?�? P  �   �0�0�0�0 11�1�1�1�1�1�1�1�1�1.2i2o2�2�2�2�233,393M3X3�3�3�3�344(4O4d4y4�4�4�4�4�4�5�6�6�67~7-8�89�9::(:::�:�:;;(;:;�;�;�;8<]<u<�<�<�<==�=W>g>�>�>�>�>?^?j?r?�?�?�? `  �   Q0�0�01I1�1�1�12X3�3�3+4[4i4v4�4�4�4�4�4�4�4�455)5D5Q5_5f5x5�6I7�7�7878�8�8�8�9�9�9':9:K:s:�:�:;;;d;u;~;�;�;�;�;�;�;<!<:<D<L<t<~<�<�<�<�<3=D=Y=g=�=�=�=�=>(>@>H>S>^>>�>�>�>�>�>�>   p  �   O0W0b0�0�0�0�0�0/1@1�1�1�1282�2�2R3d3�;�;�;�;�;�;�;�;�;�;<<$<k<~<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ===#= �     (0,000111 �      0000                                                                                                                                                                                                                                                                                                                                                                                                    �un5      ` �0  �   H  �
   `  �   �  �    �un5       h ��  �    �un5          �  �    �un5       r ��  �� ��  �    �un5       � ��  �    �un5                 �un5                �un5           0      �un5           @      �un5         P  ��   �          �� �          ��            �� �           L�             D L L  D L L 1  D V C L A L  P A C K A G E I N F O  M A I N I C O N   MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ^B*        � �� �         p�      �    H                                                       �  L    �  �   �                      �  �	                                                                                  CODE    ��      �                    `DATA    �    �      �              @  �BSS     �   �       �                 �.idata  �   �      �              @  �.edata  L    �      �              @  P.reloc  �	   �   
   �              @  P.rsrc       �      �              @  P                    �              @  P                                                                                                                                                                                                        �%��H ���%��H ���%��H ���%��H ���%��H ���%�H ���%��H ���% �H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%�H ���%�H ���%�H ���%��H ���%��H ��S�ļ�
   T�����D$,t�\$0�Ã�D[Ë��%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ��SV�еH �> u:hD  j �����ȅ�u3�^[á̵H ��̵H 3ҋ���D����B��du���^[Ð� �@Ë�SV���������u3�^[Ë�P�V�P���X�B��^[ËP��
�Q�еH ��еH �SVWUQ��$��] �$���P�V�;��SS;�u�������C��CF�F;Cu�������CF��;�uË֋��V�����u3��Z]_^[�SVWU����؋��2�C;�rp��J��k;�wb;�u�BC�B)C�{ uH���9����?�΋zϋ�k;�u){�*�
J�$�{{+��|$+��s�ԋ��������u3�����;�u�3�YZ]_^[ÐSVW�ڋ���   }�   �����  ��  ���sjh    Vj ��������;��t#�ӸԵH �l�����uh �  j �P�����3��_^[ÐSVWU�ً���C   jh    h   U�������;��u����  ��  ���sjh    VU������; t#�ӸԵH �������uh �  j �P�b���3��]_^[ÐSVWU���L$�$�D$����3҉T$��$ŉD$�ԵH �Q�;�s;�wF��C;D$w;;t$s�t$��C;D$v�D$h �  j V�������u
���H    �������߁�ԵH u��D$3҉�|$ t�D$�T$��D$+D$�T$�B��]_^[�SVWU���L$�$�Ћ�� ���$���  �� ����T$�D$�(�D$+ŋT$�B�5ԵH �<�^�~�;�v��;|$v�|$;�vjh   +�WS�&�����u
�D$3҉�
�6��ԵH u���]_^[Ë�SVWUQ�؋���  �� ����4$���� ����$���+$�A�5ԵH �8�^�~�;$s�$;�s��;�vh @  +�WS������u
���H    �6��ԵH u�Z]_^[Í@ SVWU��������H ���?  �� ����] �3;{,�΋׋C�����> tP�FC�F)C�{ u>��������5�;�uɋ֋�������> t!�̋֋�������<$ u��̋V�����3��YZ]_^[Ë�SVWU���$�����H ���?  �� ����] ��;�t;su�;suW;{��   �L$��+S�CC������|$ t3�L$�T$���]����|$ u��L$�T$�D$�%����$3҉�   �L$�׋������|$ t4�L$�T$�������|$ �f����L$�T$�D$������$3҉�H�k;�u:;{5�$�׋��q����$�8 t(�$�@C�$�@)C�{ u��������$3҉��]_^[ÐSVW�����$���?  �� ����4$��� ���;�s[�ϋ�+Ӌ������L$�׸�H �]����\$��t�L$�T$���&����D$�D$�D$�D$�|$ t�T$��H �����3����_^[�U��3�Uh>H d�2d�"h��H �9����=5�H  t
h��H �.����ԵH ������H ������H �x���h�  j �������H �=�H  t/�   ��H 3ɉL��@=  u���H �@� � �H ���H 3�ZYYd�hEH �=5�H  t
h��H ������  �堬�H ]�U��S�=��H  ��   3�Uh"H d�2d�"�=5�H  t
h��H �f������H  ��H P�4���3���H �ԵH �h �  j �CP�%������ԵH u�ԵH ������H ������H �u����̵H ��t��̵H P������̵H ��u�3�ZYYd�h)H �=5�H  t
h��H �����h��H �������-  ��[]�S; �H u	�P� �H �P�H��   8;�u��y������H 3҉T���$��y������H �T�� ��P[Ë ��P[Í@ ��H ��J;�rJ;�r����H u����H    3ҋ�ÐS�ʃ����|�  ����  [Ã�|�ʁ�  ���[����H �Ѓ�����������H ��  Ë���|����������Ã�|
�ʁ�  �� ��SV�Ѓ���ʁ�  ���  �t
���H    �ځ����+Ë�3������t
���H    �t �Ѓ��r+�;pt
���H    ����ދ�^[Í@ SVW��3���   �t%����؋�u����X����F�؃#���_^[�SVWU�������$ �������؅���   �k��C�Ѝ7+у���+���+Ń�}�L$��+S׋��������L$�׃��F�����l$��t4��+֋��c�����D$�SS;�s
�7+������T$�������$�$��]_^[Í@ SVW����߉s��ƃ��p��   7�օ�y������H �D���u��H �\��[��:��C���Z�,�� <  |�֋��������u� �H � �H ��C���Z_^[Í@ �=�H  ~@�=�H }���H    �+��H ����H ���H ������3���H 3���H Ë�SVW������<$���������L$�׸�H �����\$��u3��R�;�s
����)G�G��t$;�s�����G�G;�u���   ������o���H �G��H ���_^[Í@ S����؋ԍC�D����<$ t���W�����u3���YZ[ÐSV�����؋̍V�������<$ t���&�����u3���YZ^[Í@ 3҅�y����=   ��H �T���u@=  u���SVWU�� �H ��H ���H ;s��   ��C;�~{�s�[;s���B;t��c��   �������؅�uN��������u3��   ;u �)u �} }u 3��E ��H 5�H �փ�������H ��5��H �L�������S��+ƃ�|��֒�T������;u�C���ƃ ��Ëփ�������H ��5��H ]_^[�U����SVW�؀=��H  u	�������t�����~
3��E��T  3�Uh�H d�1d�!�=5�H  t
h��H � ����������}�   ��   ��   �Å�y������H �T���ty���Ã ��B;�u�Å�y������H 3��|���&�˅�y�����=�H �D��
�M��M��A�M���ƋR������E����H ����H �  �   ;�H J)�H �=�H }�H 3���H ��H �H �Ӄ�����E����H ����H �M  �2�������E�3�ZYYd�h�H �=5�H  t
h��H �������_  ��E�_^[YY]Í@ U��QSVW��3����H �=��H  u�f�����u���H    �E�   �a  3�Uh�!H d�1d�!�=5�H  t
h��H ����������u���H 	   ��   ���H ��%�����)��H ��tE�ƃ��P��|��  �t���H 
   �   ��+�;Pt���H 
   �   ڋ��T����������Ë�;=�H u,)�H �H �=�H  <  ~����3��E���
  �   ���t�������}���H    �7��)�ǃx t�8 t�x}���H    ��P�������Ӌ��'������H �E�3�ZYYd�h�!H �=5�H  t
h��H �W�����	  ��E�_^[Y]Ë�SVWU�����������}�   ����} �������ǋ�;�u��  ;���   ��+։$;�H u8�$)�H �$�H �=�H �L  �$�H �$)�H ���3  ���u�ËP$������<$|��ދ$����Ã�������   ����   ��+ǉD$;�H ug��H ;D$|S�D$)�H �D$�H �=�H }��H �H 5�H 3���H ��+���H �E %  ���u ��   �>�������uM�ӋH�$�$;L$}$�ڋ$)D$�,�����D$)$�<$|��Ƌ$�n����:4$��ރ#��.��   �t!%���Ë؋T$���������t	�������3����+���H �E %  ���u �YZ]_^[Ë�U��QSVW��؀=��H  u�������u
3��E��   3�Uh5$H d�2d�"�=5�H  t
h��H �����֋��������t�]��6���������Ã�� %�����;�}�ƅ�t�׋ˑ�B  ��������}�3�ZYYd�h<$H �=5�H  t
h��H ������  ��E�_^[Y]Í@ S��~�$�H �؅�u���   �3ۋ�[�S��t�(�H �؅�t��   �3ۋ�[Ë��t2��tP���,�H Y	�t�ð�   ����(�H 	�u�ð�p   ��tP���$�H Y	�t�Í@ ��H �E  �SV��؀��=�H  t
�֋���H ��u��  ��   ���w
3��Ê�0�H 3��Ë�����^[Ë����$�����S���  ��   [�VW�Ɖ׉�9�wt/��x*�����_^Ít1��|9���x�����������_^�SVWU����S�����؊��t< v�;"u�{"u����3���C<"u1S�`������S�V�����+��؊��t<"u�; tS�9������S�/�����+��؊< w��Ƌ���  �ߋ>3��Q<"u8S�������S�����;�v��7CF;�w����t<"u�; tS��������S�����;�v��7CF;�w��< w���]_^[Ë�SVW�������ڋ����
  ��uh  �D$Pj �����ȋԋ��  ��������Ӌ����������t�; tN���  _^[Ë�SV��3�f�Cf=��r/f=��w)f%��f=��u���S����u���S$����t���'������8�H t
�g   ������^[Ë�W�ǈ͉���f�ȉ���x	�у��_ÐSVW��P��tl1�1ۿ����F�� t�� ��-tb��+t_��$t_��xtZ��XtU��0u�F��xtH��XtC��t ���t-��0��	w%9�w!���؊F��u���t	��}T�	F���~KxI[)��G�ŊF뜿����F��t߀�ar�� ��0��	v����wЀ�
9�w���؊F��u���u��Y1��2_^[Í@ �%��H ��S3�j �������uj�����% �  =   t=   u���[ÐU������H �E��E�Pjj h�(H h  ��������uM3�Uh�(H d�0d� �E�   �E�P�E�Pj j h)H �E�P�����3�ZYYd�h�(H �E�P������  ��f��H f%��f�U�f��?f�f��H ��]� SOFTWARE\Borland\Delphi\RTL FPUMaskValue    ���-�H Ë���t���Q�À=�H vj j j h�����H Ð�=�H  tPPRTjj h�����H ��XÍ@ Tjj h�����H ��XÍ@ �=�H vPS�����Í@ ��t�A�9�t�9�u��AA����Ë��=�H vPRQ�����QTjj h�����H YYZXÐ�=�H vRTjj h�����H Z�PR�=�H vTjj h�����H ZXË��D$�@   �  �8����P�Htn��������H ����   �҅���   �T$�L$�9���t7������=�H  v)�=�H  w �L$PQ������ X��   �D$�H�0�D$�H�=�H v�=�H  wP�D$RQP�D����� YZXtp�HS1�VWUd�SPRQ�T$(j Ph +H R��H �|$(��  ��    ��    �o�_�G,+H ���f������#   �  ��    ���    �A������   Ë��D$�T$�@   t�J�B�+H SVWU�j���F�����]_^[�   Ë��D$0�@�+H �0  ��    �
��    �B�`��8���t�B�k����r���1���d�Y��]_^[�   Í@ ��  ��    �
��    �B�1���Z�d$,1�Yd�X]��������1ҋL$�D$��d���� Ë�U��U�=�  �,t\=�  �tW-  �t\-�   t=HtN�`q��?��r6t0�R=�  �t=-�  �t.HtHt$�:-�  �t/��=t&�,���*���&���"������������������
��������%�   �R����]� �D$�@   ��   �=�H  w�D$P�,����� tq�D$��%����T$j Ph-H R��H �\$�;����S�Ct��H ����������҅�������S�������H ��t�ыL$��   �Q�$��  1�Í@ 1ҍE�d�
d���@�,H �h�$�H Í@ 1ҡ$�H ��td�
9�u� d�Ë	���t9u�� ��U��SVW� �H �G��tH�_�p3�Uh�-H d�2d�"��~K�_�D���t�Ѕ��3�ZYYd���-����������������_^[]ÐU��SVW�(�H ��tK�03ۋx3�UhV.H d�2d�";�~��C�,�H ��t��;��3�ZYYd��������P����'����v���_^[]ÐQVW� �H �}Ĺ   �@�H �<�H �-4�H �8�H �(�H �0�H �Mĉ �H 1Ƀ} u��,�H �H ��H �H ��H �����E@�H�H HY��D�H t<}��Q�L$��t�E�U��Y�E<|���=�H  u�$�H �=�H �EH�!  ������ �SVW�T�H �� �H �ÿ
   �����03�����û
   �����I��u۱��H �Ѓ���t�H 3ۊو��I��u�_^[Ë�1�� �H ���@� �H �_�o�w�w �7�   �_^�� Ë�Q�=4�H  tWf�=�H ��u�=�H  v��H � �H j �D$PjhT�H j������P����j �D$PjhL0H j������P�����ZÀ=�H  uj hL�H hT�H j �����Z� ����   
  SVWU� �H � �H �0�H �{( u�? t���3҉���Ճ? u�=�H  t�����2���3���H �{(u
�> u3��C�����{(v�> t!�C��t��  �S�B;Bt
��tP�f��������{(u�S$�{( t�����; u�=�H  t��H �P�!����V�����   �^�v���]_^[ã �H ����Ð��H �����Ë��t�     �J�I|��J�u
P�B�����XÐSV�É֋��t�    �J�I|��J�u�B��������Nu�^[Ð��t$�J�APR�B��\   ��XR�H�����ZX���B����t�J�I|��J�u�B�����Ð��t
�J�A~��B����t�J�I|��J�u�B��h���Í@ ��~$P��
���P�3���Zf�D�  ��Z�P��@�   �1�ÐSVW�É։ω���������ǅ�t	���������������;_^[Ë�R��   �����ZÐ1Ʌ�t!R:
t:Jt:Jt:Jt����BBB��Z)�����Í@ WPQ��1��u��X�X_�y���Å�t�@�Å�t?��������SVW�É֋y��V��9�t�  ���N����X���_^[���  �����Å�ta�������;t\;tPQ�u���ZX����SVW�Ӊ�P�C�F�������ǉ؋K����������N�S������X����t�O��/���_^[É��$������I����SVWRP��1��L���t9u�ϋA�J�1��L���t	A�9�u1�Ju��t�$�w��,  �<$�77K��9���P�ƋD����t
�H���j���Ku�ZX��u��t�J�����Z_^[X�$���Ë�SVW�Ɖ�9���   ��th��tk�F��W�)�w�R��t&��9�uXJt�N�_9�uK����Ju������Z��t"��8�uAJt8�u:Jt��  � ��  � 9�u'��#�W�)���F�)��Z8�u8�u����8�u8�_^[Ë���t
�P�B~��@�Ð��t� ��4H Ë��t8�J�It2S�ËB��)�����P�H��b���X�H�I|��H�u�@��i����[��Í@ ����Ë�����Ë�S��t-�X���t&J|9�})Ӆ�|9�D$������1������D$�����[� �SVW�É։��������t0�J�N|*9�}&��~")�9�~��)��������؋R�)��L   _^[Å�t@��t1SVW�Ɖ׋O�W�V�Jx�F)�~�u��VW���_^t����Z1��1��Z��)�_^[Í@ SVW�É�1���~H���t#�x�u����	P���y���X����p�� �(��������ǋ��t���H�9�|��������������;_^[Ë��������U����SVW�E�� �H �E��}� t93�Uh�6H d�0d� �]��E��S3�ZYYd��
�����G����E�� �E��}� u�_^[YY]Ë���H ���H Ë�U��Q�E�3�Uh$7H d�2d�"�E��@�t���3�ZYYd�h+7H �E�;�H u�E�� ��H ���H ��t�;U�u	�U����� ��u���+�����Y]Ë�U����S3҉U�3�Uh�7H d�2d�"j�U�Rh  P������E��U��   �5����E��U�������؃}� t3�3�ZYYd�h�7H �E��������������[��]�U��3�Uh�7H d�0d� ���H u#�8�H ������H �����гH ������l���3�ZYYd�h�7H ��a�����]Ð�-��H ��   ��H ��H H ��H H �6�H � �H L6H �������t���������f�<�H ��f��H ��f�ԳH ��������,�H �*����(�H ����%   �=   �t-����%�   f��v���H    � ������������H ������u������H ������ �H Ð�%0�H ���%,�H ���%(�H ���%$�H ���% �H ���%�H ��Pj@�����Í@ �   Ë�S������؅�t6�=��H �u
��   �������������u��   ������P���H P����[ø   ��t�z������H �������H P�u����\�H Í@ �   ��t�=��H �t���H P�O�����tP�-���ø   ��t������=��H �t���H P����Ð�L�H ���H ��u&d�,   ����%������H P�������tá\�H �P�������t�ø��H ����Ð���H �}u*PR�L�H �M�P�H �J�B    �B    �����ZX�5T�H ���H ����Ë�U��3�Uh�:H d�0d� �X�H 3�ZYYd�h�:H ��������]Ë��-X�H �U��3�Uh�:H d�0d� �`�H 3�ZYYd�h�:H �������]Ë��-`�H ��%H�H ���%D�H ���%@�H ���%<�H ���%8�H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%��H ���%|�H ���%x�H ���%t�H ���%p�H ���%l�H ���%h�H ���%d�H ���%`�H ���%\�H ���%X�H ���%T�H ���%P�H ���%��H ���%��H ��U��3�Uh<H d�0d� �d�H 3�ZYYd�h$<H ��2�����]Ë��-d�H Ã��3ɉ$�L$Q�L$Qj h?  j j j RP�����$YZ�Q3ɉ$Th?  j RP�o����$ZË����ǹ����2������)ȉ�ÐU��QSV�M��u�����؋������PVjj �E�PS�6���S����^[Y]� �U����SV3ۉ]��M��u3�Uh�=H d�1d�!�E�   �g������E��   �E��U�������E�P�E�P�E�Pj �E�PS�������ua�}�t�}�u#�E������:����ЍE������ƋU��B����*�}� v�E��U�< u�M�E��U��t����ƋU�����S�L����������S�=���3�ZYYd�h�=H �E������������^[��]� U��3�Uh�=H d�0d� �h�H 3�ZYYd�h�=H ��r�����]Ë��-h�H É��ǹ����2��G���ÐSV��؋���������   ��^[Í@ WV�Ɖ׹����2���щ��։ʉ����у��^_�WV�׉ƹ����1���щ�1��F��W�)�^_Ë�U��QSV��E��E��)���3�Uh�>H d�0d� �E��#����؃�|�E��D�<\t</t
<:tK��}�V�˺   �E��S���3�ZYYd�h�>H �E��f�����t�����^[Y]ÐSV��؋������P������P������P������Pjh   �������^[�SVW�����������؃�|(�D�</t<\t<:uW�S������������K��}؋ǋ��.���_^[Ë�SVW�������>����؋ǋ��c����֋7��t�<ar<zw, �BFK��u�_^[Ë����ǹ����2������)ȉ�ÐWVS�Ɖ׉�2���t�uA)ˉ��։������ك�󤪉�[^_Í@ SV��؋Ƌ��m���^[Ë�U����SVW3ɉM����3�Uh�@H d�0d� ��u�ƺ�@H �\����g����������E��}� u�ۋ��������t3�ù
   ������ù
   ����؍E��W0������U�����{�����ù}� u��ƺ�@H �c���3�ZYYd�h�@H �E������������_^[YY]�   ����   0   ����   -   U��Ĵ���S�؍�����P������P�P������t4P�=���������u%�E�P������P�����E�P�E�P�E�P������u�E������E�[��]�S�؋�����@��[�SVW�ڋ���������w?�Ӂ��   ��@w2j h�   jj ��%�   ������H P����H P������P�]���_^[ÐQj RP�����ÐSVWQ�����j �D$PWVS������u�$�����$Z_^[�P�
���ÐSVW�ً���SWSVj h   �������_^[�SVW�����������؃�|�|�.uW�����Ӌ�������K��}�������_^[Ë�U����SVW3ۉ]��]��U��E�3�UhCH d�0d� ��������   �]�����
s�E�3ҊӃ�0������U����[�����E�3ҊӃ�@��	�����U�����;����m�Ou��}� t �   ��80u�ƹ   �   �e���Ou�3�ZYYd�hCH �E�   �T�����>�����_^[��]ÐU��3�UhECH d�0d� �l�H 3�ZYYd�hLCH ��
�����]Ë��-l�H �U��QSVW�E��E��>���3�Uh4DH d�0d� 3�UhDH d�0d� �x�H ������t!�   �x�H �����ع   3ҋ�������
3�ZYYd��_���u
3�ZYYd��P�u�hLDH hXDH �E��   �����E������P�E������Ћ�Y�����������3�ZYYd��
���������3�ZYYd�h;DH �E������������_^[Y]�   ����      ����   
   U�������SVW3ۉ������������]�M��U��؋u�E������E�����������3�Uh�EH d�0d� �������Ӹ   �  ���$  �׋���  ���@�   ��������   �  �����������U�������������EH ��  �������E��������t*�}� t�U��E�������t�}� t#�U��E�������u�ƍ�   �  �G�����׋��T  ���@���e���S����3�ZYYd�h�EH �������   ������E��   ������������_^[��]�  ����   ����    U��3�QQQQ3�UhzFH d�0d� �U���FH ��   �U��p�H �����U���FH ��   �u��5p�H �U���FH �   �u��x�H �   �N����U�FH �   �U�|�H �p�H �����t�H �p�H ��FH ����3�ZYYd�h�FH �E�   ��������������]�   ����   ��  ����   ú����� ����   ����    ����   ��������    ����   r   U����SVW3ɉM���E��E�����3�Uh^GH d�0d� ���<����E���������~.�E�   �E��U��\��À�E���0����U�������E�Nu�3�ZYYd�heGH �E�������E��������������_^[��]�U��3�Uh�GH d�0d� ���H u(�|�H �����x�H �����t�H �����p�H ����3�ZYYd�h�GH �������]�U��SVW3�UhHH d�0d� �-��H s'3�Uh�GH d�0d� �����3�ZYYd��
�%��������3�ZYYd�hHH ��9�����_^[]Ë�U��3�QQQQQQQS3�Uh�IH d�0d� �=��H  �&  h�IH �������H �=��H  �
  �U���IH �_����E��;���P���H P��������H �U���IH �9����E�����P���H P��������H �U��JH �����E������P���H P�������H �U� JH ������E������P���H P�}������H �U�8JH ������E�����P���H P�W������H �U�PJH �����E��}���P���H P�1������H �U�hJH �{����E��W���P���H P�������H �=��H  t	�=��H  u3���3�ZYYd�h�IH �E�   �������������[��]� kernel32.dll    ����   ����������������������    ����   ������������  ����   �����������   ����   �����峲�����   ����   �����峲����    ����   �����䳲�����   ����   �����䳲����    SV���������tVS���H ^[�3�^[ÐSV���������tVS���H ^[�3�^[ÐSV����a�����tVS���H ^[�3�^[ÐU��3�Uh�JH d�0d� ���H 3�ZYYd�hKH ��R�����]Ë��-��H �U��3�Uh5KH d�0d� ���H 3�ZYYd�h<KH �������]Ë��-��H �U�칖   j j Iu�QSVW3�UhOH d�0d� 3��U� OH �\����������DOH �L�����������H �	�E��f���������3������������������������������H �0�������TOH ������������������   ���������������؍�|������g�����|����4�����tS������x������E�����x�����������  ���H �p����ЍE�������t���P�E��W�����B���   �E�������t���P��p����dOH �I�����p���X�Q�����u9�E�������B���E��   ������l����tOH ������l����E�������=��H  uS��h�����OH �������h��������P��d�����OH �������d�������P�~���P�X������=��H ����  j j S�E��{���Pj ���H ��`�����������`���3�������؃���o  j �E�Ph  ������PS�-���S�o����E�Ƅ���� �U��������R�����\���P�E�����P�E���������׸  �Y�������\����E��-�����   ��P���3�������P�����T����q�����T�����H �0��L����dOH ������L�����X����   �J�����X���������j j S���H �n���Pj ���H ������3ɺD   �����ǅ����   fǅ���� ������P������Pj j j@j j j Sj �v�����t<�E�����P�E��	���P�׸  �Y�����������P�/���������P�#����   3�ZYYd�hOH ��L����   �m����E�   �`�����J����ۋ�_^[��]�  ����   ��������������������������  ����   ����    ����   ����    ����   ����    ����   ����    ����   ������������������  ����
   �����ή���  U��3�QQQQ3�Uh>PH d�0d� �U��LPH �$����E�U�������U����H �������H ������ЍE��t����E��T����=��H  t�E�Pj j hHKH j j �����3�ZYYd�hEPH �E�   �'�����������]�    .................................... .................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................... C    U��3�Uh�TH d�0d� ���H u
���H �a���3�ZYYd�h�TH ��b�����]Ë��-��H �U�������S3ۉ������������������������������������]��M��E��j���3�Uh�VH d�0d� h   ������P�#����������M���VH ����������������E�P�   �   �E������E��   �   �����E���VH �T�����   �U��E��'  �} ��   �������WH ������������U������؅���   �K�E��   �U����������WH ������������U������؅���   ������P��I�   �E�������������U�� ����؃}� uS��H � ��%]  �������(WH �_���������P��������H � ��%]  �t���������X� ����������?  �3�ZYYd�h�VH �������   �����E��   ������w����ۋ�[��]� ����   s:  ����   0   ����   ������  ����   ������� ����   ����    U���\���SVW����E��E��]���3�Uh�WH d�0d� ��l���Ph  �ĶH j jj���H �؃��u3��H�E��.���P�ضH ��`���fǅ\��� V��H f��^���j��\���PS���H ��u���3�3�ZYYd�h�WH �E��a�����o�������_^[��]�P��H �ԶH Ë�U��QS�U��؋E�����3�UhSXH d�0d� j�E�����P�E�����PS�ܶH ��3�ZYYd�hZXH �E����������������[Y]�S���������$ j h   �T$RP��H �Ӌ��k�����  [Í@ SVWU��0�����h   ��$�  P�������������$   Ph  �ĶH j@��$�  P�ȶH h   ��$�  P������$�  P�̶H ��t7�p3����u�7�жH �������C�<���u��ԶH h   �D$P�I������  ]_^[Ë�U���h���SVW�U��E��E��J���3�Uh�YH d�0d� ��h���Ph  �ĶH �E������E��*���P�̶H ��t)�p3����u�7�жH �U��@���C�<���u��ԶH 3�ZYYd�h�YH �E��i�����w�����_^[��]Ë�U��   j j Iu�QSV��E��E�����3�Uh�[H d�0d� ���$����E�P�   �   �E�������E�U��/����E�P�U��[H �����U�X�����+  �E�P�����   �E������U���[H � ����؅�t"�E�P�����ӋE������E������������U���[H ������؅�u�E��U������P   �@�E�P��I�   �E��7����E�P�S�����E��#����E܍U��P����؃}� t�P   �U؋E��,����E؍M��������t_h�[H �u�h \H h\H h�\H h�\H h<]H �u�hL]H hX]H �EԺ
   �����UԋE������֋E��������<:  �E��h���3�ZYYd�h�[H �EԺ   ������E��   �����������^[��]�   ����   ���к�� ����   /   ����   :   ����   GET     ����    HTTP/1.0
 �����   Accept: image/gif, image/x-xbitmap, image/jpeg, image/pjpeg, application/x-shockwave-flash, application/vnd.ms-powerpoint, application/vnd.ms-excel, application/msword, */*
  ����   Accept-Language: zh-cn
    ����@   User-Agent: Mozilla/4.0 (compatible; MSIE 6.0; Windows NT 5.0)
    ����   Host:   ����   
  ����    Proxy-Connection: Keep-Alive

    U��3�Uh�]H d�0d� ���H 3�ZYYd�h�]H �������]Ë�U��   j j Iu�QS3�Uh�_H d�0d� �-��H ��  �U���_H ������E������P�����؍U���_H ������E�����PS�g�����H �U���_H �����E�����PS�F�����H �U��_H �����E��l���PS�%������H �U��_H �o����E��K���PS������H �U�`H �N����E��*���PS������ȶH �U�`H �-����E��	���PS������ĶH �U�0`H �����E������PS�����ԶH �UܸD`H ������E������PS�����ضH �UظX`H ������E�����PS�_����ܶH �UԸh`H �����E�����PS�>������H �Uиx`H �����E��d���PS�����̶H �U̸�`H �g����E��C���PS������жH 3�ZYYd�h�_H �E̺   ������������[��]�����   ����볲���� ����   ����������� ����   �����   ����   ������  ����   ����    ����   ����������� ����
   ����������  ����
   ����������  ����	   ���������   ����   ����    ����   ������� ����   �������������   ����	   ���������   U�������SVW3�������������3�Uh0bH d�0d� 3�UhbH d�0d� �U��@�H �*  ���  �@�H -d  �8�  ��   �@�H -h  �8F  ��   �   �@�H �"  ����   ��������   �@�H �����������������   �J����������������HbH �����������E4  �������&����ء@�H ��;un�P�H ������������tZ��|U��
P�������P�H �b����= �H  t� �H Pj ����h�rH h N  jj �	���� �H �3��@�H �3��@�H 3�ZYYd��
���������3�ZYYd�h7bH �������   �5����������_^[��]�  ����   w:  U��SVW�}�]�u��uR��  t��  uB�׋��t  �=��H  u0�=P�H  u'�=P�H  u�=�H  uhdlH j2jj �D�����H WSV���H �@P��H _^[]� ��U�������SVW3�������������3�Uh&dH d�0d� 3�Uh�cH d�0d� �U��8�H ��'  ����   �   �8�H �  ����   ��������   �8�H �|����������Y����ء8�H ��;��   �P�H �������������t�������������   �����������������<dH �c����������2  �= �H  t� �H Pj �&���h�rH h N  jj ����� �H ��|���������P�H �,���3�ZYYd��
�%��������3�ZYYd�h-dH �������   �?�����)�����_^[��]�����   pin2:   SV��3Ɋ��u��t&�&���r��u��� r��9v��t	A���   u�3ҋ�^[�SVWU����$�D$ 3�3��΁�  �yI���AIu�<0 tN��tS�H�0��u��tF�$�8 �D$�8���r��t/�$�\0�9G�$�0�9G��� r�$�,;�M GF���   u��D$YZ]_^[Í@ U��ĠSVW3��E��E��E��E��E�3�UhSgH d�0d� �=8�H  t
������  �=�H  ��  �|�H �   �������  ��H �=�H  ��  3�Uh'gH d�2d�"�E�P������E؉E��E� �lgH �0  �V  �E�3ɺ   �l���j�E�P�E�P��H P�4�H �E����8  �}�   �+  �E��}�   �   �}���   �E�=  � ��   3�Uh�fH d�2d�"�]���������   �SecP�֋���  �����   �P+�غpgH �   ��������uz�ð  �8�H h�gH �U��8�H �~����u�h�gH �U��E��k����u�h�gH �U��E��X����u�h�gH �U��E��E����u��E��   �����E���.  ������E�����K���3�ZYYd��
�+���������E�E��E��}� u�E�;E������3�ZYYd��
�����������H  3�ZYYd�hZgH �E��   ������������_^[��]�   ����   a3  SecPasswordDlg  ����   a4: ����       U��ĠSVW3��E��E��E��E��E�3�UhjH d�0d� �=@�H  t
������  �=�H  �  �x�H |�H �   �������  ��H �=�H  ��  3�Uh�iH d�2d�"�E�P�b����E؉E��E� �jH �-  �|  �E�3ɺ   ����j�E�P�E�P��H P�4�H �E����^  �}�   �Q  �E��}�   �&  �}��  �E�=   �  3�Uh�iH d�2d�"�]���������p  ��  �֋��o  �����   �P+�؋Ã��8T  ��   �Ã��8��   �Ã��8F  ��   �C�8�  uz��d  �@�H h(jH �U��@�H ������u�h4jH �U��E������u�h4jH �U��E������u�h4jH �U��E������u��E��   ������E��1,  �����E�����%���3�ZYYd��
�{����.����E�E��E��}� u�E�;E��r���3�ZYYd��
�L����������H  3�ZYYd�h
jH �E��   �b�����L�����_^[��]�   ����   w1  ����   f1: ����       S���t�H �
%  ����   �=P�H  ��   �=P�H  ��   �=L�H  u	�=P�H  t	�=8�H  t�����=8�H  t�P�H ������r�P�H �������v�\  �=P�H  t,�=d�H |��H � t�G  �=d�H |�����d�H [ÐU��3�QQQQSV��3�Uh�kH d�0d� �=_�H  ��   �|�H h�kH �U��������u�U��F������u��E��   �/����E��k*  �=_�H  t�x�H |�H ��~�������=��H  u���H �E�Pj j hX�H j j ����3�ZYYd�h�kH �E�   �����靿����^[��]� ����   x   U��j j S��3�UhIlH d�0d� �=_�H  tA�M�����W����M��E��`lH ������E��)  �x�H �x�H |�H ��~3��
���3�ZYYd�hPlH �E��   �����������[YY]�   ����   k:  U����S�=]�H  ��   �=��H  uZ�=��H  u
�Y%  �   ��)  ���H �=��H  ��   ���H �l�H +��H �����H ���H ����H �P���H j�E�P���H P������]���Du�E�P��Sj���H P�������t*�]�H ���H ���H ����H �P��H Pj ����[��]� ��WS	�t�ǉÉȉ���A�� t
��)؃�[_ø����[_ÐU��3�QQQQQQQS3�UhunH d�0d� �U��T�H ������E�������K��|!�E��|�\u�S�E����������K��u��P�H  �U���nH ������M�E��U������E������Ph   hP�H h�nH �U�nH ������E�����P�U츸nH �����E�����P�@����E�P�H �   �^����M�E��nH �����E��b'  3�ZYYd�h|nH �E�   �������ڼ����[��]�   ����
   ���������      ����
   ����������  ����   ������  ����   s1: S���H ���H Pj �	�����@��tP��H �3҉P��@��tP��H �3҉P��@��tP��H �3҉P[Ë�U��3�QQQQQSV���3�Uh�oH d�0d� �U�� pH �����E�P�ù'  3���U������U���Y�����ù'  3�����6�ùd   3���U��q����u�U�pH �-����u��ùd   3���U��I����u�ƺ   ����3�ZYYd�h�oH �E�   �|�����f�����^[��]�  ����   mV  ����   A=  U��ĠSVW3��E��E��E��E��E�3�UhcrH d�0d� �=<�H  t
��  ��  �=�H  ��  ��H �=�H  ��  3�Uh7rH d�2d�"�E�P�����E؉E��E� �|rH �%%  �  �E�3ɺ   腶��j�E�P�E�P��H P�4�H �E����a  �}�   �T  �E��}�   �)  �}��  3�UhrH d�2d�"�]���0�u���0��0f����֋���  �����   �P+�؋�H�8���   �Ã��8���   �{ ��   �C f�8��   �C f�8� ��   �Ã�(�   �������tw��(�<�H h�rH �U��<�H �n����u�h�rH �U��E��[����u�h�rH �U��E��H����u�h�rH �U��E��5����u��E��   �����E���#  �<  �E��������3�ZYYd��
�����ι���E�E��E��}� u�E�;E��o���3�ZYYd��
����蟹����H  3�ZYYd�hjrH �E��   �����������_^[��]�   ����   R1  ����   f1  ����       U�� �H Pj �@���3�� �H ���H ����3��@�H ��/	  ]� �@ ��l����$�   T�����|$u3����Ĕ   ÐWS	�t�ǉ�f�ȉ���A�f��� t
��)؃�[_ø����[_�;�|��ÐU��3�QQQQSVW�P�H 3�UhOtH d�0d� �? ��   �<�H �U����  ����   �   �; ��   �{& ��   �{Hr|�{Hrv�? t�`tH ���c������ �����w`�ǋ��N����dtH ���B����C&�������w>�S&���+����dtH �������U�3��CH�����E������Ћ�������hN�d����E��׹   脾���M��E��ptH �ؾ���E��!  3�ZYYd�hVtH �E�   ������ �����_^[��]�   ,   -   ����   r:  <	w	%�   ��0�%�   ��7Ë�U����SVW3ɉM�M�M����E��E������3�Uh�uH d�0d� ���~����E�����������   �   �E��|� u�Ǻ�uH �ѽ���   �E��|��s�E��D��<_w
����uH s�E��U��T��:����U���落���S�E��D��Ѓ��U����E��7h�uH �E������ЍE�������u�E������ЍE������u�Ǻ   ����CN�L���3�ZYYd�h�uH �E�   轻���E�葻���韵����_^[��]�  ����   +   �g������������   %   U��j j j SVW�ډE��E�諾��3�Uh~vH d�0d� ���.����E�螼������~C�   �E��U��T2��,����U���肼���E��|0�
u�U���vH �����U���a���FOu�3�ZYYd�h�vH �E��   ������Ѵ����_^[��]�����   ���    SQ���$�   �Ë$�7���T���W���P�����Ë$����Z[�U��3�QQQQ�E��E��Ƚ��3�Uh�wH d�0d� �E��U�R�����u`�u��U��E�@���`��� �����u�hxH �5L�H �L�H �   �D����E�@���`��� �'  3���Сl�H ������l�H �y�U��xH �i����U�E�莼��u8�u��U��E�@���`��� �����u�hxH �5L�H �L�H �   �ʻ���'��H � t�5L�H �u�hxH �L�H �   衻��3�ZYYd�h�wH �E�   �s�����]������]�   ����   
  ����   =pWS    U��ĈSVW3��E��E��E��E��E��E��E��E��E��E�3�Uh�{H d�0d� �=L�H  �&  �=�H  �  ��H �=�H  ��  3�Uhu{H d�2d�"�U���{H �8����E�P������EЉE��E� ��{H �  �  �E�3ɺ   �c���j�E�P�E�P��H P�4�H �E����}  �}�   �p  �E��}�   �E  �}��;  �E�=  � �-  3�UhF{H d�2d�"�]���0����0���  ����֋�����������  �P+�؍{�׋Ã�$���������  �Ǻ   ���������  �E��'����ЋÃ�$������tD���  �8���  ���  �Ã�$�  �������g  ���  �   �g������O  ��$�]�h�{H �U��E������u�h�{H �U��E�������u�h�{H �U��E�������u�h�{H �U��E�������u�h�{H �U��E������u��E��
   �!����E��]  �L�H �׶��U�U��E������E��O���Y�E��  �.�U���0�E�������u2U�E��U��˷���E�����Y�E��  �E��8 t�E�E���P;E�w��E��L�H ��{H �&����E���  �=L�H  u�L�H ��{H 薶���.�= �H  t� �H Pj �����h�rH h N  jj ������ �H �E��������3�ZYYd��
�ݮ��萰���E�E��E�}� u�E�;E��S���3�ZYYd��
鮮���a�����H  3�ZYYd�h�{H �E��	   �ĵ���E�蘵���馯����_^[��]� ����   RxWS    ����   Eu1 ����   e1: ����       ����   e2: U��	   j j Iu�SV��3�UhH d�0d� �E��s����E��s����u�hH �u�h$H ��H �   �0����=P�H  u���H �P�P�H ����h�H �E�P�H �   �&����E�   �   茸���=�H  u��H �0H �������q  �E��P�H �   �������H �x t&�E������؃�|C�   �E��*����D0�*FKu�U�@H ������u�E�P�H �   菵���u�hPH �U�\H �����u��EܺP�H �   �e����u�hPH �UظlH �����u��u�E��   �����=P�H  t:�u�hPH �UԸ|H �S����uԍEкP�H �   �
����uЍE��   �ҵ���=P�H  t:�u�hPH �U̸�H �����u̍EȺP�H �   �Ǵ���uȍE��   菵���=L�H  t+�u�hPH �Uĸ�H ������u��5L�H �E��   �[����=P�H  t:�u�hPH �U���H �����u��E��P�H �   �P����u��E��   �����u�h�H �u�hPH �U���H �W����u��u�hPH h�H hPH �E��	   �ٴ���=��H  t���H �U������#���H �U��в���E�Pj j h��H j j �>���3�ZYYd�h	H �E��   �p����E��   �c�����M�����^[��]� ����   (   ����   )   ����   sender  ����   ������ ����   
  ����   ����   ����   ����   ����   ���    ����   =GI+�   ����   NoF7�   ����	   NoF7C\Bk�   ����   


I P : ����   ;zFwC{� ����   v e U��   j j Iu�3�UhڃH d�0d� 3��d�H ���H 3��h�H �P�H  ���H ���H  3����H 3���H �]�H  3��p�H ���H  h�H �<����,�H ���H ������U��@�H �\����E��8���P�,�H P������H ���H �����U��\�H �,����E�����P�,�H P輺��� �H �U��x�H �����E�����P�,�H P薺����H h��H 觺���0�H �U𸠄H ������E�譳��P�0�H P�a����4�H �U츸�H �����E�至��P�0�H P�;����$�H �U�ԄH �����E��a���P�0�H P�����(�H �=�H  �J  �=�H  �=  �= �H  �0  �=$�H  �#  ��H  3��x�H 3��t�H 3��|�H 3�� �H �P�H  �P�H  3��l�H �P�H  �Q�H  �P�H  �P�H  ���H  �P�H  �L�H �8����`�H  ���H �'��������\�H 3��D�H 3��H�H 3��@�H 3��<�H 3��8�H ��H � �f���Pj j�L����P�H �=P�H  �Q  j j j j�P�H P�������H �=��H  �,  ���H �8�  �E�P�U��H �"����E�P襸�����H Y�����U�T�H ������UܡT�H �@����UܸX�H 觮���Uظ�H ������UءX�H �������_�H �UԸ�H �����UԡX�H 辻�����^�H ���H ��]   u���H ǀ]     ��H  �=_�H  t�����Pj h   �(�H ��H �5X�H h4�H �U̡�H �x����u�h@�H �Uȡ�H � �a����uȍEк   ������E���  3�ZYYd�h�H �EȺ   苭����u������]�   user32.dll  ����;   ........................................................... ����   ������������������� ����   �����������������   ����   ��������������  kernel32.dll    ����   ��������������  ����   ������������������  ����   ����������� ����   ����    ����   .dat    ����   ����������� ����   �������Ů���    ����   ,   ����       U��j S�]3�Uh��H d�0d� ��un���H ��]  u`���H ��!]  ��"^�H u5�=�H  u@���H ��!]  
r2�U���H �,����U��X�H �3�����u���H ǀ]     ������EP�EPS���H �@P��H ��3�ZYYd�h�H �E��D�����R�������[Y]� ����   �������Ү���    U��3�QQQQQSV���H 3�Uh��H d�0d� ��8��  ��H �`�H �ǀ%]  �����  �U詷���ƀ   �E����  �  �����U���H ������؅���   �E�P�E���  �  �۫���E�˃��   �A����E��٫���؃�|W�E��D�</t<\uC�S�E������S����U��H �¿���M�E��U������E�萭���Ћ  �����K��u���@ ��U�Ph(�H h�  j
j 蒴�����H �	  �U讶����x uj �P�H P�D�H Pj� �H ��B��x uj �P�H P�<�H Pj� �H ��B��x uj �P�H P�LbH Pj� �H ��B3�ZYYd�h��H �E�   �o�����Y�����^[��]�    ����   ?   ����
   �������  U��j 3�Uh��H d�0d� ���H ��   t-�E����H ��  �P  �>����E��������H ƀ   3�ZYYd�h��H �E�赨����â����Y]� U��   j j Iu�QS3�Uh��H d�0d� �U��ĊH �����E����H �������H �d����E�P�E���H ��  �  觩���E�   �   �����E�؊H ����u`�E���H ��  �  �m����u�U�E��K����u�h�H �U��H �6����u�j �Uܡ�H �$����u܍E��   � ����4�U؋E��_����E�P�Eԋ��H ��  �  ������UԍE�Y�V������H ��	   ��   ���H ��)]  ;l�H ��   ���H ��-]   tj�M��H ��H ����h��H �EЋ��H ��	  �  舨���uЍŰE��f����u�h�H �Uȡ�H �Q����u��u��Uġ�H �>����učE��   ����j �M��H ��H �����j�M��H ��H �v����   3�ZYYd�h��H �Eĺ   軦���饠�����[��]�   ����   �������    ����   0   ����	   &subject=   ����   0   SV����؋�3ɺ   ����j�D$PS踰���D$���t�|$w3�����^[Í@ U�������SVW3҉�������������������3�Uh�H d�0d� 3�Uh��H d�0d� �U��D�H �q������X  �D�H ��U����X������?  ������3ҋ��������u3�ZYYd��3  �P�H �������l�����u�P�H ���\�������   ������詳������   ��虳������   3��t�H �������P�H �����P�H ������h4�H �������P�H �   �K���������h@�H �������P�H �   �+����������������   �����������&	  �= �H  t� �H Pj �<���h�rH h N  jj �1���� �H �%�P�H �ز����r�P�H �ɲ����s3��t�H 3�ZYYd��
�.�������3�ZYYd�h$�H �������   �H�����2�����_^[��]� ����   u   ����    p  V�P�H 3�����*u�< u�B�< u�� ^�U�������SVW3��������������������]43�Uh�H d�0d� ���%  �U����M������  �=��H  �  ��������蟤���������ܤ�����=��H  t����   ����   ����   �� ��   �=��H  t���H  3��������������ű��������������� �H 迤���������l  �U��D�H ������ti�D�H �8�U���������tT������3ҋ��������tA��������貯����u��|	���H �"�����������H  ��|
�P�H �v���3�ZYYd�h�H �������   �}�����g�����_^[��]�  ����   pa: WS	�t�ǉÈȉ�A�� t��)�H[_ø����[_Ë�WV�׉Ƹ   	�t1��	�u�O�:N�t1�^_�U��ĠSVW3��E��E��E��E��E�3�Uh��H d�0d� �=��H  �  �=D�H  �	  �=�H  ��  ��H �=�H  ��  3�Uh��H d�2d�"3��D�H 3��H�H �E�P谫���E؉E��E� �̑H ��  �}  �E�3ɺ   �0���j�E�P�E�P��H P�4�H �E����_  �}�   �R  �E��}�   �'  �}��  �E�=   �  3�Uh[�H d�2d�"�]���������   ������֋����������   �P+�؍C�8������   �C�8'  ��   �C$�8���   �C<�8��   �CL�8�   uu�è   �D�H hؑH �U��D�H �����u�h�H �U��E������u�h�H �U��E������u�h�H �U��E��ݮ���u��E��   �=����E��y  �E�����$���3�ZYYd��
�Ș���{����E�E��E��}� u�E�;E��q���3�ZYYd��
陘���L�����H  3�ZYYd�h��H �E��   诟���陙����_^[��]�����   g1  ����   f1: ����       U��ĔSVW3��E��E��E��E��E�3�Uh�H d�0d� �=�H  ��  ��H �=�H  ��  �h�H �=h�H ��  �E�P�;����ẺE��E� �4�H �[  �E�   �8�H � �E��r  �E�3ɺ   誔��j�E�P�E�P��H P�4�H �E����T  �E��}�   �D  �}�   �  �E���t	��@�  3�Uh֓H d�2d�"�]����u���+u����M��֋����������   �P+�؋���8�H ;��   �8�H �M������������   ��hH�H �U����輬���u�hT�H �U��E�詬���u�hT�H �U��E�薬���u�hT�H �U��E�胬���u��E��   �����E��  �E��0;H +ƃ��E�E��E�C���H �E��C�)���3�ZYYd��
�M���� ����E�E��E��}� u�E�;E��|�����H  3�ZYYd�h$�H �E��   �H�����2�����_^[��]� ����   k1  � E�  ����   k2: ����       U��3�QQQQSV���H 3�Uh�H d�0d� ���%]  ���te���   tZ�E����  �  ������E�P�U���W����U�X�����E��U��#����U�,�H �����E��U��à����tj �@���h0u  �Φ���3�3�ZYYd�h�H �E�   �T�����>������^[��]�   ����   ������ټ������  U��SVW�u�}�]����"_�H tJ��   �tB�֋��c����=��H  u0�=P�H  u'�=P�H  u�=�H  uhdlH j2jj �S�����H VWS���H �@P��H _^[]� �U����SVW3҉U��E��E��Ӟ��3�UhI�H d�0d� 3�Uh$�H d�0d� �E��`�H �U������E�诞���С��H   ����3�ZYYd��
�����貕��3�ZYYd�hP�H �E��   �����������_^[YY]� ����   
  U��ĘSVW3��E��E��E��E��E�3�Uhs�H d�0d� 3��E��=��H  ��  �=�H  ��  ��H �=�H  ��  �E�P������EЉE��E� ���H ������E�   ���H � �E��M  �E�3ɺ   �/���j�E�P�E�P��H P�4�H �E����/  �}�   �"  �E��}�   ��   �E���t	��@��   3�Uh,�H d�2d�"�]����u���+u����M�֋����������   �P+�؋���H ;��   ���H �M���������tn]�K�]�h��H �U��E��C����u�hȘH �U��E��0����u�hȘH �U��E������u�hȘH �U��E��
����u��E��   �j����E������E��C�N���3�ZYYd��
�����誓���E�E��E�}� u�E�;E��������H  3�ZYYd�hz�H �E��   ������ܒ����E�_^[��]�����   fc1 ������3��:_^��3�]�J[�    ����   fc2:    ����       U��SVW3�Uhj�H d�0d� ��H ut3�Uh�H d�0d� ���H P�Ǣ���P�H P����3�ZYYd��
����������X�H �����T�H �����L�H �������H �������H ������H ����3�ZYYd�hq�H �������_^[]Ë�U��SVW3�UhʙH d�0d� �-�H s'3�Uh��H d�0d� �@���3�ZYYd��
�q����$���3�ZYYd�hљH �酑����_^[]Ë�U��3�Uh��H d�0d� 3�ZYYd�h��H ��X�����]�   �H �:H `:H �7H �7H �:H �:H (<H �;H PCH  CH �=H �=H KH �JH �GH lGH @KH KH �TH �TH �]H |]H x�H ̘H     ؙH U���ĸ �H 蘟���˕���@                                                                                                                                                                                                                                                                                                                                                                                                 �@ 2�� �@  �@  �@         tH  H �#H  ��������������������� ��@ Error ��Runtime error     at 00000000 ��0123456789ABCDEF����                        �9H T9H 9H �9H    �   @   �                    t� g$X4��!rРH |�H p�H ��H                                                                                                                                                                                                                                                                                         ��  ��              v�  ��              ��  �              ��  �              H�  8�              ��  P�              ��  ��                      ��  ��  �  .�  J�  X�  h�  t�  ��  ��  ��  ��  ��  ��  ��  �  �   �  ,�  H�  T�  f�      ��  ��  ��      ��  ��  ��      ��  
�  �  "�  .�  :�      V�  h�  |�  ��  ��      ��  ��  ��  ��  ��  �  �   �  4�  D�  T�  d�  t�  ��  ��  ��  ��  ��  ��  �  �  .�  F�  T�  b�  p�  ��  ��  ��  ��      ��  ��      kernel32.dll    DeleteCriticalSection   LeaveCriticalSection    EnterCriticalSection    InitializeCriticalSection   VirtualFree   VirtualAlloc    LocalFree   LocalAlloc    GetVersion    GetCurrentThreadId    GetThreadLocale   GetStartupInfoA   GetModuleFileNameA    GetLocaleInfoA    GetCommandLineA   FreeLibrary   ExitProcess   WriteFile   UnhandledExceptionFilter    RtlUnwind   RaiseException    GetStdHandle  user32.dll    GetKeyboardType   MessageBoxA   CharNextA advapi32.dll    RegQueryValueExA    RegOpenKeyExA   RegCloseKey kernel32.dll    TlsSetValue   TlsGetValue   TlsFree   TlsAlloc    LocalFree   LocalAlloc  advapi32.dll    RegSetValueExA    RegQueryValueExA    RegOpenKeyExA   RegCreateKeyExA   RegCloseKey kernel32.dll    WriteFile   VirtualQuery    VirtualProtect    UnmapViewOfFile   Sleep   SetFilePointer    ReadFile    OpenFileMappingA    MapViewOfFile   LoadLibraryA    GetVersionExA   GetSystemInfo   GetSystemDirectoryA   GetProcAddress    GetPrivateProfileStringA    GetModuleHandleA    GetCurrentProcessId   GetComputerNameA    FindFirstFileA    FindClose   FileTimeToLocalFileTime   FileTimeToDosDateTime   ExitThread    ExitProcess   DeleteFileA   CreateThread    CreateProcessA    CreateFileA   CompareStringA    CloseHandle user32.dll    SetTimer    KillTimer                                                                                                                                                                                                                                                                                                         <�           (�  0�  8�  �n  $�  F�  I�     ztDLL.dll k1 k2                                                                                                                                                                                                                                                                                                                                                                                                                                                           0
000"0*020:0B0J0R0Z0b0j0r0z0�0�0�0�0�0�0�0�0�0�0�0�0 1(1�1�1�2V3�3�3�3t4�4�4-595T5�567r7�7�7�7�7�7�7�7�7�7�7888&8,848F8R8a8m8u8�8�8�8�8�8�8�8�8�8�8�8 9999/9:9[9s9�9�9�9�9:W:w:�:�;�;�;<<'<0<;<D<K<Z<a<�<�<�<i=�=�=�=�=>>>b>k>�>�>�>�>�>?2?\?e?u?}?�?�?�?�?�?�?�?�?�?�?      00(0@0L0T0k0z0�0�0�0�0�0�0�0,1P1n1~1�1�1�1�1222$2u2|2�2�2�2�2�2�2�2�2h3�3�3�3�34#4+4O4o4�4�4�4�4�4�457&8e8u8�8�8�8�8�8%9:9N9V9l9�9�9�9�9�9:::O:|:�:�:�:�:�:;k;�;�<=
="=D=x=�=�=�=�=>*>>>t>�>�>�>�>�>�>�>�>�>�>�>�>�>�>??!?<?D?p?{?�?�?�?�?�?�?�?�?   0    0'01060U0Z0_0�0�0�01)161�4a6r6�6�6�6�6�6�67@7�7�7�7�7�7�7�7�788888"8)8-8G8P8Y8e8o8�8�8�8�8�8�8�8�8�8�89H9c9m9x9�9�9�9�9�9�9�9�9::':1:O:T:g:s:�:�:�:�:�:�:�:�:�:�:�:�:;
;;;";*;2;:;B;J;R;Z;b;j;r;z;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<*<�<�=�=�=�=�=�>�>   @  �   0/0�0�0�1�1m2�2'333@3R3n3|3�3�3�3�3'4�45�5�5�5�5�5666.6;6A6K6Q6V6h6�6I7s77�7�7�7�7�7�7�7�7858A8M8W8]8l88�8�8�8�8�8�8�8�8�8�899"9*9=9H9P9c9n9t9}9�9�:�:�:�:�:�:
;;#;0;B;_;o;;�;�;�;?<�<�<�<�< =$=B=>>A>O>�>�?�?�?�? P  �   00,0�4�4�4�4�4B5g5�5�5
6Y6l6�6�6O7g7s7�7�7�7�7�7�7878F8|8�8�8�89$9b9z9�9�9�9�9:E:w:�:*;2;7;<;A;F;N;S;�;�=�=�=�=�=�=�=>>3>;>T>\>u>}>�>�>�>�>�>�>�>??"?;?C?\?d?}?�?   `  8  �0�0�0�0�0171c1�1�1�1�1�1�1�1�1�12z2�2�2�2�2�2�2�2�2�233;3R3b3�3�3�3�3�3�3425>5Q5]5s5z5�5�5�5�56X6t6y6�6�6�6�637A7�7�7�7�7�7�78818Y8`8�8$9)919>9Q9d9�9�9=:P:]:j:s:|:�:�:�:�:�:�:�:�:�:	;;;S;[;a;s;|;�;�;�;�; <<<<7<m<z<�<�<�<�<�<�<�<�<�<�<�<�<===#=+=}=�=�=�=�=�=>>4>I>c>�>�>�>??<?J?�?�?   p    .0:0M0Z0a0p0�0�0�0�0�1�1�1�1�1�1C2Q2�2�2�2�293A3V3�3�3�3#4=4�4�45K5�56L6l6�67!7&7N7X7b7�7�7�7�7�7�7�7�7I8U8b8o8v8�8�8�8�8�8'9�9�9:%:8:`:�:�:�:�:�:;
;;*;�;�;<-<5<:<J<R<Z<d<l<�<�<�<�<�<�<===-=?=G=e=p=x=�=�=�=�=�=�=�=�=>>*>2>B>d>l>t>�>�>�>�>�>�>�>�>�? �  �  0000#0*02090?0G0M0S0]0b0o0�0�0�0�0�0�0�0�0�0�0�0�011 131>1F1Y1d1j1w1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1
222&2-242;2B2G2]2c2w2�2�2�2�2�2�2�2�2�2�233!3/343B3R3Y3o3t3z33�3�3�3�3Q5`5n5~5�5�5�5�5�5�5�5�51696P6W6�6	7L7_7}7�7�7�7�7�7�7�7�7�718<8N8k88�8�8�8�8�899E9M9_9�9�9�9�9�9�9�9�9:*:2:E:e:j:|:�:�:f;t;�;�;�;�;<&<0<<<G<\<g<�<�<�<�<�<�<�<=F=�=�=�=>><>T>b>�>�>�>�>n?z?�?�?�?�?�?�?�?�? �  �   00Z0�0�0�0�0	11�1�1222&23292X2i2�2�2�23#3<3P3c3v3�3�3�34d4l4�4�4R5k5t5}5�5�5�5�5�5�5�5�5676�6�6�6�6�6�6�677T7�7�7�7�7�7�7S8a8�8�8�8�89!9+959?9I9S9e9�9�9�9�9�9�9::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:l:w:   �      $0(0,0�0�0�0�0�0�0�0�0                                                                          �un5       
     �    �un5       �  �8  ��  �P  �    �un5           h       �un5           x   ��             ��  �            D V C L A L  P A C K A G E I N F O   &=O87��$B�:�  �       ztDLL �Uupdate  UupdateConst  �SysInit  �System  UType  �SysUtils2 KWindows UTypes �Reg �TlHelp32  �SMail  qUnitHookDll                                                                                                                                                                                    (       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                                                                                                                                                                        @    @        D@  D@        DDDDDD@     � DDDDDD@    ��LDDDC�@   ��L��K��@   �  L��K��@       L��K��@        L��K��@        DL�K�D@        DDDDDD@     � ODDD$@    ��O��B"$@   ��O��B"$@   �  O��B"$@       O��B"$@        D�B$D@        DDDDDD@         DDDDDD           DDDD                   ���Z7�Z��������e��f���j���$������o���"������ �n �" �� �� �n �" �� �� ��@��x��x��x�nx�"�� �� ���?����&=O87��$B�:�  �       Hzt GMMSystem  �System  �SysInit KWindows UTypes tUinject2000ExitProcess �OpenThread  UType �SysUtils2 �Reg  �TlHelp32  @Other  �Uconst  NUnitMain          �                                                                                                                                                                   