MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ^B*        � ��     �     ��      �   @                      �     �        @                       ��  �    p  ,6                  ~�                             ��  @                                                   CODE     `      �    PEC2O      @  �.rsrc    P   p   H   �             @  �         0   �   "   �             @  �                                                                                                                                                                                                                                                                                                                                                                                                                ���>�Fx!��0��b{2&jĥ���V�e��֍Ð��J=���ʖ^i�s�.����ג��/��,�;m��&0��y��Π˧��n�I�����_&]�u�р|��8�	/�z�~���B�:���,+��u����cr�e-!� 3�>��)lCvRi"+�rc��y���5&�3���i@J�z/J���߅��I�[���߆2:PXG|ڍ���گl�{U�ug��	1�XMTJC��9�3I�ޣJP��Lo�����A�5� �C5Pӈ�N��ٷ
\��J�}rj7��.ܩ��1#I�85�ꛣQ6E��XՋ�o�|���o��p����d�Pt@΂�NFY��8��<�i�.2�ݞ�g->_i/qV�b=� 2'ڒ�|�֝^���=��[�l�Q4qO���U��}(�8ټD���%ʨ���T��_6��j���6Єn'&;�U��k#�*�A6s���u�v$U�ʨ�Ǌ��T�����V�q��j���?x�-�1 �)�[���=�����U�d�	�4��KG?,�N,���H9�ʓ����m5��
2���+�������6������� ���@B-�E	~p٪�����M:�e,Z�3(�-QS������ilU����$n�)�R*Jq�as,.~��;�=����YS,�UJ�2��.!l:�����-vJ���1N4���9���6g�2��tm�^�{C��!�����,v�
�Vʽ`9� �I�D.�R�N;_P}��3�.�ɔ��މ���H���c1Q��8��O����g�Q,~�h?]�7����pYQ6`�J�U�=����0�K��S'̗�)ޱ Ӣ�X��8G��~��Ck��!cg[k,�0UyBa�����'��� �V�lYŨG�W�-L�8]�e�"�3�A'���o%�Zn�*z$F�Lͺ�u�CChN1Ъe����}`��޾�&79�ݡtMr�.�����T}��tˋ�(��,����Nԃ=��:m,�LTZN��t%��N�Z����������񼠵[I�]�:?���94̥��	���6H=	�+�r~�]�
�����ML��f��?��޴�D��|1_�� �O`ǃ�FҸ�Ĉ�JK�*�W�2
�N�gݷ߉Dn�C{&�fG��[�tJ�!ji�Ux��&wtTgE�}��*�g>�\�z��e�?�ٌ0G���|���7�r���Y�hu� ���8����k�J~�5Z�\�����2������ؼõ�+�]x�o1�.�s��BvP�����Wr��}K���z׏�-�kÕ"���	��_u�z1�db����[<��ӂn�+���'���a�V慎ژ'z�O5�7p�i��KsR,4���mR�v%H��5�8՛qߵ<T��0X�,���GT]O�{�a�goJ��g�c�I6}�8L�� �ɂۂ��e�ap�^�'0_Z�&�X�`'٢K�M��^-�︳'�sT����V��܃���Ѫ����et�0 �#��E?P+�c��|bD�S�XX
�ɵ�ݩ�ݫ��#,z�Nͦ������}�C}�!������0䍙뭷R)�ւ��)�!l��[KM'�Waz~($��)���n�h�\�a������-�0���W�=:"臋(,ȱd'��Jf���q}m�h�6U�.竪/���z�.�QN�qf�������kű�y3���="&��l��0fڷ��v�#�Q���8��mC:�T�y�^�8 q�0l��z�NS�&��͸`	��cv��7�}p�ja��F/�M$�c8>S���$f��UD���f4�*
�^�m��<1�GYO1	,]ɸ^��Ӄc�f	��i�?�7E�O^b��R.i�ҚH�o���N�^A��_iq��po&ݞ�Ӣ����q��Y[�g��9g��3�����u��� Fӄ�[Ï��l�jZ����-	g''�EM���jj�J�(��3t��[����,� �&��y����=�����M��j�PeSvz�vD�<.�U�bz%��<�P�Ҏ(��䝪$��B�Qry<��=
dOҷ�s*�I=���ޜ���v�Y�YzJ�X=R�~�\�n�%���� Q�0,��u�xO�&�2�}*
\���;�Ί�?~��)��H^�$I�],9��)�2�~S��y=�� n`�F������E&D��i�v�߀���d¦E�G�G_M�TD���,+�ؚ���u$������Ջ������5xUQ��ΓA�LUH;���Μ�C�>�x>V�V������H҄RoR|)�oZ��DM_�����RL��ybӉ�B� �\3��YH�&�N�D�V����;����20g��b�~V��}�*G�L��3G6�=��'�0�%�I��b�����
�ϔ�z�W��uQ[^g�rB����U��ɏH�)R���u�Q�˻�����������t��+p���'��J��M�u~��x�Ƅ�Ձ��r�T��O��g�e@O]����u6�u��SU�� ����b1E�������l�:���><K%���S�Eh���֋�@� %�^~���帾۞.5�':)/�#�Z\�&߅  ��AB�l��21��Z�t�r*q�i��c����H����܏1����vǹ	5���;O��0�O�@��65d��<b�a��] nո�T�MKV.DL�^,���~B�f�₺ti��Ӷx�����z�͹b���!�Y6���%rX�t����H��Ȭ���4�/\R208�t;�q�+ؓ��C�����*1R�+�ڃN�pe2:kB��*([�"�A��C�3$�M�U���֜�R��Ө�;�V݌G�џRP.5�Yi'I�F���5u	�Ab���&]�r>"Z@�#p�s(J&s�� �C^�l¿�5�ڃ�"�0UddJ��t+εwi�h�+K�<�!�#�r��)l��6�bC�ׄ�b�{��as�H�PX�wX; ]�qؙ�p����`ĸ�[gsn�~C�К�Xָ�`�2�z���d�Y'M��[�����~�HX��d<	q+RކuZ���܅U�ހZV��
����qZ��m.��g�q>��`;�h��Т:�x?-�� ���ZC@�y�)�?�=%���_���D2󯲗94&�/����_�����TL�������A5k��2HPU�n�����|�p�N�#����az������e��v(�ȳ�T��Cƕ���{���1�G� �⥪�uJ��Q�E�<�s��~u���Q3�y�L/�W觖`Rn�X( �' 9�S�ݷ;��
o*N�~�Oh��IZtgD�w�~BI��z
���`�h2J�E-Ŏ��?�0�9�kY�j�(O�\��@���A��G�5/r�־'�%帪��_w^��u��!6�	�0kV��h����5������ࡃZ>!� Ax�d��)��Oh8��Q�,z�A>Ě�S������,A�'���p�Tv�s���=L
������imd� )��69�#$/�9�O�-�"69�G
��:{��U>��6�.A��2� ��h��`���zW�ʈz����������Z3NTv�6#O fl��(���j�]C�lB���I����?r9�kߋǰm�4An�!��j衉����S\��oˑ�H�3�8�c��7��)d���JB�����mo�����/�<��Mx�A/���ǵz�@?	���c�9�zLlՇ�z��O��N������<k�瘍kT�(-F������t��ߩ!�~�ёo/�82F�S�W�RMV4�*]4�MS��l/��Ѻ���F��`�i�~ hu5�x5 ��yS�J������.R�$|nS���e��A/_�Ф��*��T�6�޺�-��>,�d��@��������bxk~$���}akN����y��z�ZlF"#"�t4>��ٴ7� ىy�����-%����db�~�HX�"4R{<�t��Z'�p�3	vu`�:��L������ \�ݎ'W��~(
9W�Lqn7�q����6%�/�5����n��?D���X ��$�Gg
)�4@0ur�3'��T��jf�ڵU:sL���u�T�v8�����T�g��V	(����=t�T�������ϳ-x�g��7�ޝ󦹭����6|Y&�{b�ƪ��}c�)5Zo�f�#��,�r��j�>r�y&U"j�~Rv�k�n���#r;��D>.?�r�E��g�+��M�I�:�%20A��Bt.K#+��e(`��ӊ��gt�!�IC8��Ġ���0�"����f9�"C/�RM~q8n���rm�j�@ߟ�����|��MGP�i�.�C܉���(��
V�T�{�Th�`����0�<�n���~H��y���$O�.� IKPee�G\	bI��J�}2o�Y.�(��)�}�,A�z ��<���[���g�[=����O��F���ۑH]�(�h����i�^��������7�����;���N�76�v� ��:�ȅ��a���7��*"D���E)�"ܧ�����.D�^ X
3�'m��JYTV�6%�
���v�T;���뎌A�!�{R+IE�������}�/�n"�n:�^�%�r��>#�U";w���s���w@��X��	�X�H(:�1���k�u��T�k�OT�̡y�($�;����q�*f�P�o�AȬ[o��w�:b�<^X��K�7����YC�sXk�Ɔ���M~h1�Z<��}a�$(ܘ�b>yݧ��V���w��dD�xĉﯩb�eO�J�9�Q�d諃A�զX������T�v��1;]ݐ��d�t��!�6�Sv�e ��u'��L5R����KT�Fn^�`����0�x�M��d x��A|�����p�Ϭ��1��TxV�v�K��kq��GM伷@ � ����CF��5~B�N޹����'���l+?�!̰������I������GBez��Gi��0�xpYj�`q	Jg����"���(>`�!-=2��4|���K��y`���dB�^�����=;z�@Щp&v(����-�E�����bu3��� �в0V�%N�v��y��vʶ0�e%fWSl�[Y)��|�f協ڴ>D�8;%&�-`v����G�MX��=�>�P0~�cr�}T~L����&vI�ɀ	"�ZdG���PN�z�SJƝ*Ն�Ak���TH|0w/f���D��njl��28Ë�C/�)�=�ǈ��A,f:?�u���I|{r�b���*P��R���3�+9����7�f	�VKUo��i��>��a֋h"�bƎD��폗�-sh��MlPb���I\�l8L_%��Pp�6*x��`�.��9V���K;���n�R`���]����q)c�|��q�'�B��/���G]�m��^�B��ex�ʭ��m�� �0���%���rP�b]M����������kg9yBI�tgkU#� ��gN�~��&�fW���60�7 k�)�F���a��M�3�b�8�e���ʉ ���\�.��=�3���a3H��걐=�aXl�{��CxޅP ��nm�_�0�t��S�$� X���M=ɧ�~kA�ђ@-�Rg���b��v��D�j����.t�nps�'�9�3�v�g�������1�&Ef��C@d���U�-}0�T��^ۨᮣ�ym��ص��ˉ�T�Ǫj}X�T]p=�I�[\�~��T��1b=Ec�&�N������~��-��G�S�7��K��hjC@�Tn�	#���F�{���F ;Oj�Q?K�A�Qm�1���fo�+x�݉%
sC����!c��B��.!Ã�������I"aBgn�)"ͅ��M�I�yK�Yx�I���Q3��Dށ:;�\oς�A:��\���#��QuL���:x�XA�/���J'�PFW/t�uH�+��<�vE���.���m��0�!�>-�.��]lrG'�%��g��yvHZ�>B�F�fO�a���v�ۏ�%|��~ "F`I!�5�n�beF V��� ��sa��
ӵ&Qi(h�ozy��ͻ�D<x�fX'��wp�gg�x��aoJ��f�ї�����d<P���D4)d��o�Z�+/ڀ%G${��2޸������d�'�n��cch��i��X�]�e�٣�3N��j���V_�!* `���	7Sr ��)(��[0�'%��.��ԭ���:uʍ9eq_\�� V�Ԅ,�G	!F�󆳈�B��D���%$�ry}2]�oZ�#N�R���k;H�	\�
�����5��h̵U	ѧk�<�b�����SCP}���J�d��I\:��o�Dь���$L3��K�O_�L[�jѻMgYƎ�#>���ξ�8d� ދw�iQU��<��O聃'S��Ϗ�����ErV�J q{�@�`f�5��|�f?Q�cһ�,R��W�JP�$3��<Z;��c`�kt�i:�b�]�:E�Z�֛�&u1P�eT{ȃ`�n	*.?B&�+l�`��/��?�op��l�-�pD�t��H�/`�D2�(�( �#�� ��iB�9Fӛ�Ց�Q����f��6b�Ԧ'�~\Tn���*�����p���G!P�`+'y@�]��`n�I�Ke��ʛ.�[����3�) s��}t%�(���4��~	5��sp~Fp�XL_t&ڭ����o��}�;���5RҰf}kQ�.Cc=��ߑ��y��F�%���To���32o٩���ph��U��ᗙF��==��U/5j�����@��꧖h"r\|�,R+�}i��W4?j�
nml���Z�u���b �!�(��+��e�>�����.L�� �q׹�U��B=�.(�s	�87̍av7���qo>�5�z`J&�.@��-ӝ�Ӂd�Ƌ���[���b�4��:
��,��0jQ��C��S��ܼKݒÿ��h����><8Ǥ6~��#�ϩ��;h�*4�	d@V�É��wqc��h�;??C�����a�x+�5���S*1f�I�.a������D�c��"
�(c�=��I�`)-��+��~��9G_�<���^���ڥ��/9���mef/�l�B�X�)�bע�?*����N�]�F�'�;G ⴏj��*����t'����z�2>�nN3j��H�Pmk� ���_��y�+��+��Բ�:D1�`����ƾ��ѫ�X�{:�l��(��8�2�b*�S4��	������Ջ�ա�{�s#e_S����Q>C������y�[^�~D�I�_���oQDM�S������_y�� P�4x"k1]�<)�[�X<X�z��ێ>GK�r(�!��_*THE��dژ��	Z�g�g�q�)�X׮T��S�nx�� ��k��,!�;�F�0�t�L�{��Z���G��p�3�<�NxZ��":`!#��z%����(�XWUc���Y����Kf3��� �0�H	��O#������e�l�����?vu]1�n��Y���:����Z�&<l 'L��՗�n�J���k8��f�U:ȃY��;�"AZ��/U9j[A窩�Ѐ:�]Z��1���f�`G�Ug���Pd����K�/.��jP�e �aC�� �tD�� ��]!�
���UgNg�[W��)���BJM�a2��'�M����VCL
�n�ab
.}I�׸сƋ��_�{�r�L�C{ۯ�4��v���oL�O3�?lg�$
p����֙�$h���ސ7�D��s����!�`��� �:��4����֫�W/FH���f6�dWZ�	�V5/K>1U~t)�B/�`�$�Ə*)����Qik�bAM_�un�q ��yb��]sk	�B�M���Y8�s!x��O���fG� �#%���.�~���ר��/�}�)f!N�ezK��$w��c�Χ)0C{E*��e����z������h3)��A`�E�)|/��Fz�O6�g�t�XD�D���������t��C����g���=s����X������7��$�#e��&f�|���71��`}[x%n�Ij�wk�Xѣ�|��*#����UP]���7s������&	��Ō1֫vI:ץ��`��$h�|a����1� tn;�	@7v�V1,��"�,K��}1��[���:�:����f��Х�n�B�LwŌb�.f��E�@K�����*����������fI�޾��3}-�Z0��lJ�����\	���=���g�W�޴^�~���� P�u.��V�x�_i��a�a�n�5�t(���ɖ*�o8���+,�)���]$΍�ju�c �,��ё���v�X���k[:�4��*4�*�#z�fٙ{J)@�%>���7���[�1Cx�E��{�o��O__bx;��t��A8��L�!#7Њ$���\v@�
3�a|uQ�D����7�g���lW��/�t O[���4���g/8� F��B���
Q*�b.��X؀�� ��zV��MjZ�z6�#\���*M�Qk����:1a=IȤs�~���_�9��	�����O��vb(n���\�Kur�6��%1)�<Ɏ]+�ƒ�j<;Qc�^��v`��P�Xj��o�pS��}��'��������F)��2=�KF�2���P��{�{=��s�Y�X��/�&�(�ߐ�9�b��u	������nP�&���ld��a�BY3Ȕ'���C):� �y%Ԣ��e|�>���eF-���Yv6�G�[k�KO8s�� ��KU`���)L��do��tťu:ce~����S����;GMǥO|�+��{Ÿ�p!KW�rѤ�������4�/�6��V�E���݉X�Ez����.V�(BHS|��l���n�*���d�Y��� f�Zc�ϟ%��%�*(\g��)wG&���<���&����q���,e�̬��o���W��]4dhN�?��E{XBa�LA[A�Co�0��S*�h��>�:�*}3�S �v'��hJԳ}���p�?
s���8��.ɰ��P��k�>�B�}B{���:�����X���g����\�~�EX;��'�����/��:aU��
�ׅi3鋃wD�Qk����W�
�����03����;1$q̑��"L1�Av������,�=��A	w�B(�g��"�:S|�U���D�>꒳(Z3�ۧ�}�m�:X��*l��4�d��й���g����;�����9��X���n#4eL�n9G�I?ñ߯�}�<~蹱,e��r"m+��2��؏���X?��������W�f��-d�I�(5=��y�}�3R;�1I`{ū7p�mHU�c����B�*^l���g�'ܥG���s���*8	�v�����|���oM"��Z�eV��Oc��Ǯ�T/�c�(E���(y��J+Kó`��|ua��5c����%v� =�P�Kx�����b)���������k����(�׀�6nKה �ƋK�{Pg�~�����Z�%��yd�@��ɺ���=o����c\j_����@}���C���`�[��'C�j&Ho��[��J�I6>.&������6=��-�Fʃ��
�!�{�"��I�|�$�ni�]zB��9�����(z�^L����!1�@p����ȣ�J۴(�!.�χ+�����h�¼����<�R��ۃO(ۚ;���j���ԗ\�����f���ȶcn_�)����� ��妫�^��6��ļ��T��:J������Z�D��ѓ��ǴM�H:7�b�֧f��[M�5��>�hV!�����K�a����#�w��X�|�o�\[�/�lI���}<��?�ɗG@ �}"�6xc�}�W 6nƶ��#l��@�	���C��XO������7�����.��b(��j.Y�J�v����S4ٗ�)��Ya���DT��"�$RA0���>0B�B�H��t?j�C�'��I�Ǝ'`�l�Nk4��1��H7�U
Q�e�M���FKѦ�~u������t��o�0�|̻�6z;OX��6^m�H~�S X�\����_���xq�_����6t������+�#�]�W��!��� �NgO��1-l�w�+U�	a�̰āїc����ǘ^&��t� Ib�]B4�-ny�47��ԏ�h%(�xK𓖘 `�=u��VW�K�V �˵�����
B��c�0xUm���=<x�kÚ��pDw]E�s9tn���LR��M����e�5�5��:��G�o��)�h���@qz|��g������jK�K��]#�',4b����TPt�y�8����m�U�R�]�7-��#�{��
�{�}ƨ(m��E9� T�*�#�ˆ���n�G�UD\)�[�q,��9�4m����g��H�9
�hp���ϐ�5���ܮ��?��5���5�(�avL�o�7��O����*��--��["\��oq�H%��|q��%X�V/{ӂ�d��'�\Z@r����9���߲�]��T~�� pGz!�(��&�U����4C�����^'��m��<}hP�%�5&��g�j�
 !��l=�<��vl�X"Wr�ъ�:��E?٣L��>�g x��0��b�?�����Աgh��p�������N��C�l�/�c�{u�#�V���� �x9`�,���+9.�<���;�P�?|>^
�P���s7��B՗ZiC)'ͺ��X��6��@D�����ә��"�ɿ���F�+��B�2�u��6�-�&�'�!4���]6���D$Hr���b���=�-[���) ���2E�Y���-t��l�߻�C�~�c����k�8)Ԧ ��ԿzH>��ʏԈ�����	8k�|k��1�y^�.3�#s�>r^�;�MU�
,1�}�p�lYi��|��������Ñ �����H�fV|}pה��u�$F�h�ۓ�Vм�$�󰤥��sG�K�썃J��o?�w���-���w��H]8q�U��j	$?e8k�@���DA�ռ�,(Ef,Rw�0gQ(]�&�ۖ�i�
�!�)v.)mՐv��|�F��ê�@��n��\~�m�E_3�pvy�]���B $��z��{�|�w�S�]��r	0�K�TǛ��y�ݯwP��|d��}G� �
�2,R�ב�S>�햿|{>)��uLe�%G��l�X`9ɳol�QCZ�֢����n?�q�z�*�U��#b�8d����V����a�~�k^��D��EgC�����6�;6�����O�!e��a#Ȭ-~m�a�Ƽ���?@��ITI�)��0�O7/�\.4� ������n:[�f�nH��6�~K{�fx�����,i2�
�{���˃�p�S��"G�$�A5>|���H럠���QΫ�Yy#�p'ږ���Ѷ"� �v����,��᳉�V��wBh/,@�0�'/��t�қ�M���F7�6f[��N8
Q_{���!ݾ�M(�7�ܫ?��J�7$��D�$Q%p2z���B-�ݑ������_���xύ�TS��(REv��t�QxۢR�(�M�"5Ŏr��w	�Y�5�>�kL��R�f �wOػJT��j���,

9C��+"˼��B�/g��IGFw�$C���v�C��͙������'���L�Ϡ ��_�>Vq��>����K�y�&Z�!��W/�إ �O	6�ڛڰ��'�B+غ���f�E�[�t�ӛ �����^����3J�qyy��m�⎰dɇ�^��\�
�Íͣ������ﳾ�P�R���ݚ�Ҹ?�Oh����D@��ŗ�U��$A���Uj|"q�C���=KQ�]��n��Q�BM�B�U��H��������B�O_X�f�@%�Dh ҥ�-랩z�[�P8K�O�^Pcm����=o��	��$�
�"�������{���a80�/���6v��ƒ���@0��Y�xW_F���;�U����=��C�9q4�e"o�/+Dm�V:!�vN7��n�<g�mjE�1e\V�<�4�n��׽ک�@A�:��R��C�q$ߤ����S�A$g��G���,{2O_|�}@I]c�lEU'�W]���bf����b|�� ]Ĝ��lĺ,�P>�~�$��,hf��3�������,t�/���W:�$ËW�զp�r�mAO��0[~��ȥb%��Xg]����%d�n1� һ��\�9J�ܻ]Z��X\o�����Pp1�2=�}i�/��ְ�^����Y���� ����P�Jy�Y=�����������态�t��w�A���h{ȉ�"� ����\����-������������z��f09yF<����7���I׷��Z
��]X������@roᐋ�	S�}�Ot����<b5�C9 A��Ѝ�׋���gȜ���K���z�h#w�L4��b��L'����7��1W��g���%��쐺����Ӻ,Z�r���EGK����T��zcY�W`���<jTe��C�7cX��VP���~Ga��a:
8�x���%�}���&b�?W���ή1K�{,6?�	̭C����I�1�4%wk�ܕ!~N�+7�����;Q�5k�	�ƅ񰐘˙�},f�r��|4$�np�n��$���Ew�΍�\=��gxdޮ���J����1�$�Ѕ�X#OXO���OsZ�I�/쬏�ǧ�?�8�pI���3�
�R�m^Y�z~Y:sP�|O��`��p�2%\�����d��]�a�=\xu	�o�M��w�^��&f��My� ^�sHG��	�������g�7%c迨s"������v����Q���Ps��fB(�B�d)��aD�G���_s�>�w�u�!�n��9Z�:z��AeW��,5���i*t��O��*�d�;�G�緤^����~��1�l:z�w���qu�ȇh�z�5��m9���>�Uu����NZc�6�xс�����h�M�h�?F��\>+�%{5#,�m+lHIQ<;�h��ѵA��e̠yS��=�x��o�������DZC����������/Ҿ%����4�ك�,��G!]<��tU��ša�9p�*%�8��R���򎴾�Lo��ę��U&���š��1m�g������Ò(���=h����C�f^�Mg�C�<�~n�Xl%]\���,[�p_��^`j���@����y��0g��|���B���"�-q�\z�Rӟ������B�&�_����3�g�����%��%���X�-r���9vv��b�۔�J�1ԁ�c��"m%�*��A<z� {[���)��x����M��;�e(����1=&º@�X�,Oԫa��8+ǫ�,ȥK�]�t�s.�ĸj%���_�+t79�c'6�C�Ff'�짽����f��(}&'|P�4�ߖ��;'���g��yc)��M�\,C� ���:,���9��j@G��4K��t�51_��{��Q/J��X��~✆���k��4�G�QIH�R�N82�h����Ln�8���.�h"5!��� X8����w݄W��׸������ևEa���\�%�{뗺��J
1��W���Y6J��B5�6ݰ��g�ٔI�ɟ� P �	rp�i������wL%��JYL�+��*�;gɱ�����%L��b�Z8��>�b��,�w&g*��u���'����:�+����:��8b�z t<k��
���v��_�����Z�,2������N�����+F��v]DC�/i0�A�"U�{��G��/�W�5��募	���o���
�V�Pf4*I�vM1�T�|�m�Y9l�؀w��t�>�k�|�esW=�d6��\��>C;�t��I譲�2؆x|c2�<Ѵ�_{QQB#�KL#��mex)2��ub?�o]�#��J�������ެ#��'�r�-�w��%�h�ow)�gu_!V�g����{��Ͱ���@݄puDEOk�<Oŏ����2U�D�����f��������Mxz�cr�rG>�L���Jg�`^F��V��M��<F���JCt\W���`'ʛ9�<��rD��@
q/�*�|[|#F�zW��O�6�
h+��x�C�F��vu�mz��m)�a�-�N&�W��8 Ɖ֮��D���#Bc�x�F'�yfS~�Mv���װ���L�X��Ȉy�֑p�YG���T5vC�6|�Y�V&��R����c���\�����K�d�֛2xUW�����e�%��F,�G;{��0���D����2TV3�Lf�H�&����	c.O��T��xyԷ�%4�[�Ћ��1�v��l}�&�=<&�r�Q�"J���7�Ǳ�fuW1���k��aXP)oe�S�J�/V� ��k<������\cz~�E7$�scH_�wn�Q��>�$ YT�`�LQ�*�V���؉��ѴD��}�*���$I�k;�<Qdއ�G�SS��Z��$���ɶsF#�ט8��>Y/�3E�IF������	xf'0K��V!&0���<��	l�T�8��z��\��R��X؛ꬍ}���#�8��;�!��IZ��bz;��� c�ؼ}�PZ��3�2�D�
bS[QƵ�MT�׫i��b_~��z!�G���R������G�IJ�t_7�D
A�6�t�v�(��=Y�f"�N��T�"�Q���]�ܮTU=�
�i{�`�C��rky��)�б8\�����&&J���qL~?�3��r��0��(�,j�G�ia��`�I�����s���2Є��J@�ڐ����4e�=����,B�"�ieEv���Ax9`���ޡ�.9�۷�р��lx����!X���@of8�T�q�')�j2��I�����}l���-,[��@b5���k���X5(H'�\P��뒽�H�wϋ�1\��L��Y��łO���[��jU6ȷ�����IM�c_*cǟ�
��@;A5X�z>mBHe� 
�5j4�
���d�~��2��#�M��5��a���猦+`��	*��ݪ�.Md�ǎ^9�:�Lj��ݰ���Z�Sz9��PH�і�:;�y:q)mn������;x>l�`�5���b���z�Ϣ��Ǖb֙�ԫF�麷r��KاO.4ۼ5��""��U���LE�n����S5��)4�:���d�4��"ӆ��m}D
����:e���[h�a��$%��"��^���ףE|kx1V�q��gvU`���;AW���+Y�P��<B�Y(dx��"n �ΐ���a1�����0�<��ͦw,��§����.�� �G[��#IZ2��/��qp���{�Õ���ADk�'�M�6��LH����6�-�1��5�(R����l"4� �X��V�Ãi�g1�nh�}.�x@��ה=Bb5�q���9��e��ͧ-H�1�V	ݨ��=q#��$4m�$mO��6~n`���TC=|��s��ۉ��������b��w%�Y��� ���0D���{0��"���!$�x.��<�U�vI�����9j��bI��`8�E���F�*�Bǣ>I�V�Kq�TV��9����q'�����0�n��t�Д�&.�\�����j��1�:��J <5�&�\]9�z�6}��<l��LM ^�y/�=���|��1[�%b�e� �\(Wo�,q��Xw�-�2E�zCI��˦'l����9��K�
����Lte�m�8�o�Ji��yhL�R����[S����P���|�����/�f����c�b'?-��χ'`;��}Y�l':������h ���C
S&�(�j���qE����m��f�b�-=��LbL��*b��J\�9hu��)"5��g�[Nu��Nܧ���Z�A�8�����S�+�_6A��x) d͐z����~у�^9��2����xDjui+�ٴD�:jN����N-��K@�{���R���^�ϱ�����@є� ����^�a��W��F2��mȥ�����MT�%V�{6q;쯜������C�����b<�M�Sӿk\ʒ<�:�l�;�Ms�R�Ѽ~�]j�\��>t7Ro������}%����o�����
���2�}����N]�ށ�|�X5@,�tC��{��?��p�[g�p<�=�ZX��]����q�6=�V5��}]/�sif'f;�6T��Tv66�����e]���νJ{!�����ߓ��E�,�g������������C5J��{�yӧ����O3օ! fb�^�nR"B�Ӌcp������H��ڝ��?_�p�f6-B���z��t��k����1�������cr$N�ƅ����"S?�����!��,���P��'���u��w_o�~
�!��,����� �ػ}&�g3�7d�����H�m+LxK�ˆ�Z���0��Ra-;��^�#�^vB������vH�<x��_~�>	p��/xOC����y�&-Pj�C6��ri	�1�w��`�VH��B��4�����{e���d;��b#g>���J�]�"X�1-�˅��MǕ�u��<Wv�g���1tQ�J !P���ՏN �駍��Q��G<�3|�����uYqD���u����G�i�i�/K|���vP���m]E��v���Dq����|�س������iG:�2�^���U����0��N)�}0��E�?-�?�^�~ �!��q�8iտ�+,�z_�v��z�D.�g.��I>�&��4S8�!ٴt��������S�|�s��K~;��r�^Q�tQ�� \��Ew����s�fI�� �4�m]�Z�TW���IF���xig�`*t2��"#&�ߕ[¢��'+b�#LjB��9:&%�k��@��~m;����ӐY�R> o?⽝QJ���{u����32Z�����rӈ�6��U�v�ח\�B^�y��@�zL��Q��z�|���. �Ȍ&�J��Q��J�Hz��*P�;�H�2 ���槈����;���jTu�N0��?G����4���m��`�Y��=�P�5T��xi��s�k�Y^��a�M+9p����b��թ$�8�3��%|��&~LT>� �}�pwM��g0���	�j�V�rT�͛�8c,
|C��2���x���Z<���T�*�'+-����TK�a��Of��"[��b�e��:B6����	��r��H70�(���Xڗ��b"Z�no�J����G � K�:-*�w�foR)倪V�k<3-��=[��Y�l����s��R���X^F��Hpz�����M���S��T`�gM��d�u�u[di�\;�л�Zڴܼ�G	W�����V��tq��t�r�p��0��MW8o�
�_� m���m�&�^����y=��`Y�s��#:gm��}w�aD(+ȝ�30�@]E���d�cɔ@#95{˾C����HT��+%���$��� A��uīQl�1{0H4a��Nr�_�sB^H����O	��if!�m�k��l��Pt�	�I7�^�ϩz��ն�f^�398	�MV�,��;O3�f^��]�Ms���s�|��Us�����v�����?���A�'w�Q���`sl)�5��.���;zz(z�y*�����ޅ%���0� �jl��U�����\��cL?u^'р�������$���@�ZA�t���u$�^�EXv��q��ͤ�r$6b�x�ZC�琺��"XͱGM�R��L��h�@⫝̸�$��%\�.�y�J�0�L���~��qZv�P���QP풷B�3�̰ fx��L��#�����wJ�h��=9���O�7�x�z�*��OmCt�g���{dy�אb��((�ǂ-�4v���r�-e���Hr�m�K��w�Gz��F��J��\�l����q޽�S�;�n��5�Wd: J�0M�qž��P�˙��e��ѡ�ؤ
��O�D֋��sH����u7z�)��M%}�P8�6��� -��8�T.�؞X]��ǆ&03�Ao�H��3g>w��k��ɩ���?�(I���h�ø��7��ڎ]�j�n�(2�s� 4~�Tk��YR���#-���
F���ڲ�7H{��5i��V�`<����̞���0=����R���i?T7�/��9��M�Stn!����$P�Z�>[�9�
/r���<�(�7̏����3٧(��Х��_�"=�\h�w���D��m>���[�$Y�	P+4������]��^���2��2�Ӹ��_SE��muWl&��Tdk�Jq�>��I��q
�-���� ș궓a��II����vu����d~�r�M$��I'���ॿ]�+�$�g�ѝa��!4�dc�7���X�ϔ`u����Tj��!$a�Թ_.IFg�F( V�B}rW̫Y;�)�N�R��@��,�"��w͂}��W���,0��`[$�����x�C�����^�n�^������<���w�Sr"��lτqa�6a��PCw����M��3�����-�ZaRk�QV��Qge�iP���*z%C����wƕ3]v*����C��6�k휢����p�Gz�c����N���k���!Z�iz@�k�������*axV�î2���1!QB�S�a����F���H�x�����w��;�
�2�/��^uNW#U�-����Z��$���x>�]����k|�
�ă��� ���3O(�M�9I�O�3�O�Oɬ�d�����W�J9�B�)���b�|w(7�삔n?�z��1�aN��(.���X�"�2E���.�?�A�� �4\up^d����y�@!�R�t�Q���dI�]�\�P[��2�I�>��uD++��]�b�GR���t=�08{�V#LZѷ�a��&��	Y�y(�S�S�!ʀL�8�~B���l�����G��hDh��-�K,���@��8�r�|��a����fկ�0]��1.H�Z?S	����N��XEF�iYz���L�C��ˌ�:4�&Br����{�4��?�mW/v��ń�ݛ�O�G>-f�N�q�B2����@+,Q�f�u�$���7�5A�U>�u�\ H{2Fܞ�������W�!rKYb��;=Y���$1�kf�_���:M����@�M:"C��(�].G��L^��F%,����4Q�"������aи8Rի0w�f�;9D{l�[�ZR���?Czt�x%�ÅӐ��6�iC(�\�	m���v�kH�s��A-������Z���'O`j�v�[��F���B�5n��?H|aHt/�N[�_���q,]GۺS	�J�m���Zt�����?�$y�c�����u����<U��37�	!�XYd����Z;=�C����;Ӂ�GK0y�h�gC�X�e��������dچ�P���|�/\�O~�aE��(���oxdQc�����$�+Vu�������7���B+߄Ml�z�������O@�p$�aK�'� ���s��rv�����{w�ҢONb{�c8�}��X1���[-]y�ʿ��Y^�L&�{�e�9�$��^�7�a�]��bd��"��X5���	B���-;^W��x��;٪Sr�8B�Y�g7����L�� 8^I�Y��T̿BJ���,xVv9
�Ï�~����NX�
Ok\~ß��3J����$�ύE���������*p	����wH�l>�lP��N�
|gӎ�8����N���&xʦ�A��� ܎M�'j%�rG��鏵��N�
WYcZ����==D^zcѮH�cD���6x��N�b��d�K�Ϩꎺ?�6�������bo�&�7%���cI\M�d'�Q4��Bb����Wk9�hpd�Rl*S�e�^@;�C!���ֵ`����� ���8�v�%{�7��_̓��+����4�=��'�S��l*���[~�q�fuB p<!�����C�u�rO5,pN�M ,~n���������LO6��z�6�]��-�2Ͼw�5l���Z��DB��Ω�D:�q�$�}�BA`nG��������څ��=���徆.}��v��=�4W1Ъg���<J�àoI� _���Z6��B	,w�>nJ{�����fas^�̝)z�P�6�K%S�U��}F��f����K8=^V��U��_$��|���� *ʲX\M���9���mfzO��#��~�>W�5����U�8)�7���V�D9X�΂J2� ��b�q��P�:�O:�1LB�Ν��,�d�Kˈ�`P��ڨw'�=ʽ��j*�i�.�E���=�y���0N�"������w��j3S2#<�_dӘ����K�/����?&�u͓F�D-�S��OuU����P�a��l�}�Ə1X�,��Q�l<~���?�].�Y�k�$�vP��� ����?:���,����û�&2�>�b�2���"wx0�^��A8믮>@�QT��<��}�[d��RlN|� ~��.�6�~�eT�b��,��v���|B�v�u��`����m�qp��}~r���U��l�A��,6�1���h��8�`�8�E$�aa�w��7n���Nj0�{-��^�2�2V�ؕ�r���?���>����%��e�l�4g�C���3�s��!��"�I�@�9�p�8�sW�黮M���@���<	���n������i�.)��=�N؝8��T�S�ہr8B��e\�Zj\]/�^��F�����>w�퉬�N��B��:n.�6{�I!��
f݇O�{�u�
ZuA���(0z��5}'��x�3|SB{[yVd���/��:�W�"�]�B�ڞ�~��.�O42����I6Do�{~��l��������v�$͎J���G�}>-=�˻&bcw�x(����/z$*�H7 s
\ ��� X3�DЉ�X�A�@�׍��X���-�Ę��	�L�-��ޠ��Fε)�d���!~j�tpx {�	�^+;���-k���[�Q�#�6�տ)��]R���죶;vX�9�vl��޼�!-����7�M<4�*��2K�A��cX��Zpn7ͅQ���T�{���ܒ��V�4��A
Ɖ�u���c� 
'pCbb�܅�	��=G� .O�'
5�������xBr��R�.U��J���F�-��U0��c9���\�j8)��0"�if�� ���7Ĳ��D�/�o~T�1`9w��+��Ǥ�\�<����P���cǶ�@x`P��&�UI��S�;͜7r`2��93�k��z��.+h#�;P��V��xE9���W�n����\���URk�v
%��rV=�����28�Jl Wy�����O��-��q�N:��<���YC<b�X/�pX2?����Q>�<\^�P���Dĭ�R�߲s1�svA�<��7��qb�AD�DY��F(�!#�o��#@���'���",j���0m>'C�OUE�d�~\iLE�vG�|y�o����=3�_��^��� h_Y�ߗ��k5��� ���k���#c��Wv�"{���v������œ߈��~�Q����*���lz���'$s`ܞ~���������Q��>7�L���6�Rt1�aJρ�L^��{0㞷��u�BSe��<N,���2˨
�ڠٻ��='���@J���@�|���K��_4�U�C����xp2P��H>�����p�M����:��Iҋ�3��&1�j m�rtI��` ����}&B�k�	�`o�R������Wo�d�ǿqᔽ'Rki���`��wYeς��(�ؽJ�#��W�$�/���F��G��e��[N��Yb����@�/B��ư|.3e���<���C�>:���X�Jn�Ò��e�5ܑ����ۗs���~�[.��/�,�]���������|���9�}g��Mg
sb�`�R�#�N����q��l k�I����+�����)��6d�yF/��,�(�(�\��p}�=��pd�͠�
s/1�Аv49��_�򾖎��O�y�`廏c򽬆�eT�향C
1c�I��.=�CY��_�����њ��7e�!��ƈL���H�@��)�P�L���?d�})!�՚
�\�a.r����^7~X�´��kC ,� v=�fQ牂8���Q��*��b�p��
b��ğ�3 ��a[	ct������^%![��멘�Z��NH ��ۅ��h?�.�Wi4��k$#j�]����oK������u�	�m���U����ZR�cN��͎`�'�h1d�����+�)�iѭ\H8R�]�ca߮k����Gt���b����A�-����}�{�=���Ύ�M����`+�ܱ?�~�������>Pr�f2��LdϐG�!�>�l-�t�#[�龣�=����Ĵ���>㯻o���&$� ��&+Y�@ϡF1��T��&>���9�e�	���J�ؚ��ʏ;.�������iF�]/�/P�1��5O��|{)ҏ�c���U�p=9�V��28����1���_��e2\��v�xWtgѹ��;�~��<��1WE�Tv�^�=�RW&��T�.���,���!�e	N���Y�\�����F؀���Gݮ�!�j���u��P4!���Y*.;<��"h��G���H��{:�op�Te�@���k���k'��z
��I7H�O��]�j��"ٮa$o�~>��a\�Zo:���
j��e��Fc2�R�#5y������:)�.:������{��Q*v�r�G8���hXOd0�F����f��_h�H���'V<�уp�ƪ���]�bN�2ɐFa�L�L���{����d�q\e*��,W��<��2Gu0|�f|ew��`J}�NҠ�&!���x�	y�H�~�I@���[#�QO���p4a��iж���qB�T�C�Kl�׶ۄٚ�i�'����c��o3vސF"L�"��yb+z��بgf�x�24R@˵Y��k����N�-�&�Ͳh�b�^Vu��+�"'�3yf�ھ4$�$IW���H��gA'�:~�D^��k`�	����!O`KD��)Q�����)<�^�>�ŏ
�[ط�`�֫J�}ǗmZ���W�u0��^�Xýٵʫi}�@�D2:O���)i�Oe���AL��n.�M�Vō)�A�Bi���H�M����Ѕ��o�f�㧓��7sZ�
�(;����]t1�4��/�*��=my$�Цi <��՗"�W��������Y��jBD�,�ݱ��r3^XP�pж�bb7�k���[�Zm�t�2�Q��6�`Ex:}�j~	_U�^ �t���s�<-���%����B-�/��1�4iLi��h�B�$�y.rGt�����?���pFM|���ElVƐ�
b+}\�)��SG��l�-]b5���U���|����4�>o�% �,���@����wY�sqR�<��}rc�C���<�'�!�5�N�ݐ�Ij#��	E��U�u�]
�l��Ѳ|2��B�6c�|c Jߟ�%x��~}]U�.	��b�,8S6�1�WѴ�<g�"[�T�Ȁ�=��9in���򢱨�,�C����2�e��3>L���=ֈ�#�'�~ZFE����2E��������m'9<��+/դ;'e��t��D���¼�S��93� ���W�t���w�{�u�O!�*��s�N���N\��^�&�lA�t+�R��{��v�ep�?�\VBLj�?���.���j<
X+���x�G�XK+d���w�e�-f�Wʡ�<��$]�t�f*YP�6B8돵���Wٍ�x�����;�FB&X�^�Ԟ��H���'��#z.������ ����f��%Q^�2���q���)?(Ŗ��J���;C�8OT(>T��|�UAxЁ5&Q�T#�����d�4��_�_꜋�S�#v�k3��,������ú��Q\i�(�@��/)&>f����D�k@I@o/���׃7�N;�bc��o��
�v�yB��s0�Ł�2�d��ж1�cgF��_n���&��k��|�oDA�Ҹ���]�q�|�d�pv$�_���
�+֫"��A��nc;$k�sh���f{�!|���0�߱�Ӿ�{�Md��٧ �q��'����5Ue�	�R�10?�Ss��?�{JO$s+���&��2�0`,�,ge��?���	޻\�5M<@�lO���Q��wf h��ҷ{��g�;<z[�ݞ Ș�|���,�����M���fXJ�X	S�ѝ�`��p��ג�����V���F=�����X'���,zh��5#+��ʴI_�k�
�9ӤX6�Rg��fT�e}�#�	︀�X�����']�(��q	=�)�	�m�D)ݫ�@�Im�4�P���T|ָTFV�עM��d�ݴ�<���䚙ϲʤ�1����@�)06��%9.D5d��P�P�V��!����KT�n	����T� �+B���͹�U���9�J�#R�j�;�/FU3+�sH#nU�p�!U���@^��~(d��9$k��#����U�z�j[�	d+�o�����Ư��F���ǊUx��B=��LX�U�K�"������������#�w��>�g��Bl]*�ߙ�p�V.{?��f�m����t�*��$l�{\rP(��9�7�Ԯ��������gf�.�7�!8�lJgJ\!��,�{�A�L>����U O~2�s�̼�3��H�4�ӻ� �"&um�}8�dް	�������t��HEY�1�$�Y7�-DޱKR`�y�z �#��/����\�/��<W��C���w%��{�f=~��J	'�������J�,��PCo�AXi�A�!���RBtyd�ۚƼ�G��{�^}#�i��mi}�E�GS��L����t���?�:/���HY�T}Z�؁C:�}�w̻kC׌���{:�z;P�����U�y']W<���Շ��/�e ��sT�ej^hB
���{�����I����i*n�'I*S��j;�+W4��Tr���Gt
�����U/�i#�>&��s\Հ�����A���|GA�&@��έ,;��H���b���39�V���A�+�lQ��q׿���� 0�">����իR��ց.uz�b��6f<���8*0ƪ��ˉ��LX�hr5��^UW�M��j���n�{��_	�7Q�T��}�lOx�ˏ�hvfYی��{��M&��y��]S+H���/��+��<F	��Nl2Oxze�y�GIS�9�7��S���re�qS�� �>^)�d~&�q�v�P8����jg�v{t#��CR��/�5�37�q6:7�`gh��w�x���<�'5�0������	x�u}�����ԡO�8��1�T�"��CD�M6����̕�HԖ��(WS�DWJwń�q4R�ɭ��T�<���d<��+�|v�)�DISm���b�`�*�����D������L����,6*.#H��w���Y@��K��^���i  h� ��S?R�2j���X;}l�(�����p�r��LH�r��0x��] ��ဿ�,H�.���Nr����ds4����<Eù++���@�����M�*k8����X�7��m���d~c���?��a �Zy�n\�����oNv
���F�8e*eNv;	��.�X��Oy��E~��8h��A�΢c�׍r<Ͳ ��&'H��/���"��<`�lE>�ٛk8�^>J�E��l�~�`%����̝9P��E�5=)I����r/.mΈ�W]Q��|2x��9j�����cI�(�TY),aF���I����B�Y����O�����@IN�����'�{��?��J�e/s ݐEx�ќu"�f��g	%;V �	PO����S���g�\����w�����{>Re�!>^��T��� �T����"plͬ�;Hp�vb���݉�Z��>�X�gFO�0;�7����"���������(+���윈���m��0�<�	-�QsC��o���W����΂�fu���-]�~�q����X��i��5t�t|+����Z��:��r͍�R綒3��=ɗP���s�Z��u�v��ICfBOqą�R��Dpy�F�lv8��%��ۚ����:Pv���xw�$Y�wʁ�@@�8sT��V.�܎�!����^kY���b��J&��X08�~N�0� :<h�#m��B�3b͇�����Ў�DvJ��u�.^��Q����L�(����l�ln�p�{A|#�#��O�X�%J�������_ƺ[�}�;�T�;��G��O�6�ᠦ$_�
@I���l�9*o	���y�@����O껾{j�F�wC��?��`��Y�X5&=�Y�Y+��1�%Wb���Y�Gu�r)m,1LJ0�~�)����l��ZN�h�	�4��$&c�p^E$n������x�)K�t��ՙ�]ݣo�Q b������:?���䐏���NDT����R�Y���
���P/k
l ��5t���Ng%�`(��jI<p���:a���$wX���w��ç��Eɇ�T;x�nm.~ҕ��n�}x�C�
�+[��ѥ��q*M�����5��w��yY\�b�4;"��l�O���tEQ��1��=��coZaէ�X#��L+OD�K!�y��]�BΨ�l$qyϚ=�i�(�m
a�@��� [Y�I���\�����*�J�*e��:�^s/N����,uzo���_b�ѧtY�^UW��S��C�
#�M3$�-���1"�����r��Jd%�
��W߯G���i����'9��˝|���ex�Z��h�~9��˯��h\V;I�T�R�!7VȚ�w�Ѫ���l)b�5sM`�'�Me��!���aF�����	�ښWs�Y��p��Q�A�6�����+��%�/=�4_��wO��߰�S������h�v�ЙM���U �M�`٣���<8lD+_��Lx��E��!hEM�{w�^�7�<�t��If��HI�A��E׎73!��&ґ'[��!�� AЕ^��P,��F�vҡ�������D@��a��=��dr��I0v�>��w�<n/tEN	.@��F�/"_c6��h�J�u/��}V-�o��M��)�0{��5*>�@xʟ�A^��𬍻=���i��*��e��6?8�LA=��@0We���:EК��֟ř|�y��j�,k;�	������w6(�|�eM$�"��!���������:�b;)"����������8����<������(��[*0>븈wk��V�jw��Z�뀱�����횰�'S��l�b��H�YG���!u"'�'�����(�����lDm::�y�(��W��� g5��_�[+���QQ��:p��c��T�E��n�rxn�b������k�Q�@FA��vP����(+�j������Խ�?B`�c���d�$��Ő۪�Cؼ���5/�ڌ.3���9��U�[z	o%"��a�7Pc�FC<%9��]����>���x�-K7|{0�E��V�����R|؆���F�b]�E�ը�@r3F��J�� [}����$���$U�}j	�|9�.F	��}D�JR@��J���'��t��1<^�c
�be؞�C|��Lb�U�p;��a������ �|�K}j�z���C�Z柧k�̆ڥ�"*Z:�gʨ�l�Б�F|�h��o��� �[�:F{�X�;v46<F=���V�O�ϵ�1]��<�/��B#.��:���~�5 �D�_��-O��o.��F4���͝/2�q+c�ǿ�\10��
5�m�-3\�qa�K;����ę��,a����"��O��cO�o�9R[��߷'.A�3�! <��&���3�\�ڽb	��c�_�)��uv�D�iINa��H��䨂��2#���'�۠ə���G�Gmx��ڇO9�����?k���ғ��xպ���`��ʣ���^��0=��x]pu��v��.�aή��9ek5��x�;A��R��V�v|�P�<�X}�Y�i	S'+�o1r��܋20�S�̫���0��H��P���4l'����:��m˹+G��.���$�hi����EfZ�8,�֚x%��=��Y����~˻
|�c��ħ�^��5f:R��5_=�ǃk�����-��v[��NAN������y������S�%����N���!�������xn���2y��J2vObb���~;�q��O�z쌯jS��/#�qu&�,��n�Y�\
X8#�fo6���k(�P��X��4��Ȣr�z.a�+Ow��)yx���P�	z���: ��;*$��%�+�Kz8s�����r.cޮC0�ωJ�����q�U�H5E���[�p彑Rs�?�=�'⨆�Ҽ&�4��nA���,�D���I^���<�==����ݮl.�P�w��X��d ]v�{��6��+�����/b�j%LWBa~M��'n?.��%S7O���\I��TN�s����M��t�V�{X�SR<x����9���X�u��QsJ��������07�(+�cW�@�	�5pl�D�����A�h!>^�{q�s?�rD���]&��z}'y�C)�u���<'WH/��=9Z�ϭs���0��&�fuS�̜}�a��x�N������@��Ԃ��vH�]pUCh������ �����U�A�+�����A�d����k@�H�ˀ�%�U��j�& �K�|
$�p���啰�(G0����;��Du��ܲ��qx"j�@{���~տ�yE^6
� �с�L>�ED	��A)�$1cRt��Mݲ������$��H0�F�3���xF�*�w}��,�z�6[`��ͺ�˂N��1f�� ��!)�^��Kj��	�zGu6���E�~A45�� ���4;��j�s`�(�ߛ��OSc��uU�����D�R��g��R���Jh���|jO�y��P��Z�jK���4q��L�a��PQi��b?u��O�/No-���gMm!�U�T��r�H�;nl��&��N)�A�J�(��=̆�;�K��q3���N�*a�NJ@]"��t��}$�<.�SC���X�Ny"�{n_ŏa�n�_/�S�6��S\H@�~�@��}��C*�G����[!�X�h-U�~���6G�vV�wSv���A�9t���-�.��\3�0P�_� ؇������3O�]�Rv4�뢜X���B�!g�
꜅�'�Q5�(��EŜ��?{1�o7O�^;Ȃ���rC�J��%�C�8ݫVZ����M��O��Hi-#�1f��)��NXpZ[�'H�g�x�L�>)�����c҈�f�,7���"�����~~ۡ6���F-m�bw'D��fy��x�P�*����������'�JL��V��l�Y�E4i�,x�Qޝ�0E5g��߰��[��<�t���f��t���\U%���v���g���^���4����V�#;��[�_W 1���P�&LU=W�
eſ�" �t7�0�IƳ\�|7��H�~�
��{�T� E��5�;�|.��k
6�(�\��XA �B�̥�[�yw"���D�IE��Σ!s/��{����mR�Q>�e_�����G:5l�i���J��0v�<�,*z�v�D����)شS��Bp���e�=yޣ�:c�ErQk�a��X��p�t��+dD��b�+`�*����X�SO�Ɠ�����Gr{��(a-��S���"�!�C��� K<C�˖ ��5*H�Ȗ�����zgia���\�!��kl��3CE�e5�Y�v����\��x/�N�~zLz_9�9@�+3Z��98�X���|n����Iٖ�B���#���E֝��5��1*�uI�7}�^���Y�(+�f�� �to�o��珥�"	�S����!i��!O��7D�)�5��!��)�[����L���l�,��08��{����_98�+��^~n���u�ޢa8�S,4�7����~�q'��4�#(!�`�����DI{M�z�u�<uvںDC�I�r�4Mh�T�(��n�(�"�vg@nl���q�/��6���}k�� �� W��ԮI��n&U+���Ui×����*�\U�D���2��U�;ԍ���W��f#� F$���R��B}`��8u��y���e�[)�0�Z(��x�1�t���Br1�l�ױ������i���չ��M����0Xgr;���a�tc����n�|Έ�1D�V�:J���2%|?Y��o�x��%2�+˓�`(m�y�SƖ&Q ��,��7��+C==C�PL�W����O�ԭ�y�0R�����y�f�0��BGnQ=!�-�D�����^�H�/Lf��	j
0��I��}����~ﴞELH�fE]�홈HR��Y�D<}?65RY�D�Eg����'�3u��s��3g�_|��Y_u��1��ڊþ��l�e�����T.P��VVOv1s)�7&��~�KsΑC���'#n�y�\)g23�l�����]MV���.�WNK�#6��E֐f;��j��Mez���mw�����=���lq.� �߮*!=�sk�m�a��o�8�C#y��Fn#	���
��c�d�mϠ	�����}�Q%���c����
���ȁ�xp��O��qFn(����l��W'{\��}�+�싩��,#9d���?�����B9#�;�;��%����4�#Ȭ+RU&���б�aBei�h�[���*ۯWT�GDӯ����K�ߕ� ����}B�g\���ŽN{t�¬�,_
��(jKֱ��s���c~��zϙaP��?�>P��蜸Y�b�w�Pg]�k�1��qi����m�n�{��]�Jllp�q"C�5.����f�iߢ�����9S�Eb
�25�J�Q�LUAE.'
���E�&�A�c{H޽+ݛ�֎�����2S�'Ai$h���mT�=rSMa�DW�"@&�.��}�)L�-�`;��>U�q��C�xMO�K�c�i�V�^ݢ7��`4!-���i��\y�@K/�K_�P\B��|p~�>�h�٠WU?y�N�$$��Б�BI�H�jP���=V��j	�����ߡ�D����u�.�6a�-u�1lL�_��G��%\���e�9��V���9�f����I�zy���v?��{-����Š(?x.�}�ڿ�1��0��|{2�5�J�q:$�	{c��;o鍅3	O�l9�S����kU���sz����x(<�%'5}˞�%��ށ�]d��љ�al~�����	W7���2�*67���-Ӛ���3���u�P[
k�����Y6a��~T�K�~�{��]��E��������zO;��R��k����_D2^�?`�)e����|����{h���З������ѩb�ؾLҭバ��B?�*��c�zH�;�;I*f�dZŜ�N�dƟh�]5ǌK��v
m ^���N_ �����(�'�w�'Q��h ����cz��])�{����򱳓��-���69�.����QC��]j�mApA���Y���������5�ŉ�����w��
~v��R�0��@w�>ȱ({�c5�����Kp����EQ��&\!ț�QBZ@A�Q �6��<���"'��e���}�����DwW�|J��xm�
ťM+�r��X<^�"��n�t-��r{�ru�ͻ������jd��)�,)�<��N!�6�39'�_TDE�?Pa�Y��� +V��Y�foT	��L��H#4ЦQ���!����噼�G@��D�:�k aB��X���l�[Ei�Wr{ry?@�i�������mH��a9h�\�W�%b�����<��q��>�rgT}#�T�8n'|�_�SԆ����9��-�-����|~v�Ҳ����d��EU.p��W<�x9o��Jr��y�����;z�0D��1�f4`F�����`�����2�����c��'�Dc��#	C�� ��W�!_����������4�ZT!ܽc{���Q�ŵS��=�;�˞�к����`����}�xj<^	�鈆LGܩa�����_� $Rf������~�Q┥������i1���/^��DU3W��2ײa^���[���Ζ/���.1��ō�:���D�x������H��E1�ZV��;��k�OQv���(�V�zq��+,мSe�"̀56�M����0�~��x�<a�XW^a	m̎�m��Yqe��c�v�׍}�7���'s͆]f���i��y���}f�f)�Z�Ԛ��f-+鿢+t��<�L)��TɎ�x*�l���_�� ,}J8��\�eP���~�.�)z����9�3(���и(�zF����*�:h��6?H��r�t8�)lP �/�	��_�$��1�ȱ�!�im�>�+��N�cՑ'���J�z���3K=Q��D��GS����T]7�#��:�i�_� ���Z���[h�}�$^�e���U�P��<��Y��3D���|��ąh����$������a#��=�`q����U�~ib�%>�ϼu�7�3s'�����6�Q�(��D^��L���`�H�#��vIğ�h0��tb��4Z�>G�Z]k��j����#v)'G�S�q�q�'c`��wo�ɰ8�Y�i'��sO��9$.�z\�c�Pk�"`{p֒
�x�P���? ��4�`����$��{^�:��B�j@���1�}?6�� 
����ڃ���qs���q��p+�8r�tu61]qÚQϙ��?�^�2�7���,2�[FB��ivHy�9 "P���Y�2��CB��j���V�}a�x����
���lx�k�����[��l�?g�`�)�I�*H���B�6�*���7r;�����_�`���lݵ���9F�z5���ff�f�P�����/f��Dj����]E��[PEJ��6B�luM���_eU��?/��n��k����9}N�]�2�J�-�/� Ζ����W���cͳnv�4�)`������Vy��:rk���$���2����P�#wcy5@RxD=�_
���
��OD� ��h\R�@�oɲʥ:iR&9�B��g�u���~}�4�nU�kY��}�qz%k�zX~��,,�D�=߈�������~x���z�0�FV&���a\�`�9�"d.�iKI��|2�5C;�gR�� ��k�@�,�H���H�m٦���>qϳ c)Y��q��G�(U%�9�1��_� �}3�0��[�3��e��^�e6c�Q)�c"}�z�%G��Z7`���N���>���ު5�%�P�(ڇ%��f#��A)�)�"��=g������@n�,�j
.��a{3�oe�����E��e7ڶ��Ek5[��e9F7�K�3�GU�<�Arqi��3A�����!ƣ<vUK\��
�eD���o�:�����뷅.�KV;mUut$,"E۱�A� p1�����1f����lt2Z��r7&�鸍�E�K�������6Nr��':����y@�?-8o��ڭO�C���f/�4p�|�����Z{�}��U#�ԈbF_��W�OQx��p%�2�2��I�)u>@���+����*�,B�-��j�o>��WͩcTG��L�?:�� CW��Kf%���8�^�f����r�ػ$��;���Iq�ؒ ;٭�_�\�ݦ��Y��&�7��bW�%f�6���	i�~)4?��7���@;�U�ڎa���+�����Ǉ�uYcW�q��B��<H� �=����K�;n�y;�^��<����´������'�_be����x�{�Ap�,z�3�	!qr9�\a�<g&~oX���a����z"�GF��A��î=N���Y�N\@��$$!%�'~���Ǎ�`��U�t�㜼ǳ��7a�ᆳp�B> V�B����d��T���
��x�����<i�)�Ae�#E���NaD�r'�h��s#�[C����T	9/��z�K�0�M5"��$��F(T��U������}g��w���{S��5q�ɜ� (	E���+L9� �]!��C����Ԙ��j�V�=������A+Ҧ�2�����;��g՚$�%��6/��@���ҫ�/���iSʁ�E#�0cF;��r��=N`�/��7��5Ғ�NVS-T�t��?h:�F���7�ϣ�ģ��_':�/M:?&0�'��J�΀��ύ'����)�>~��(�S�b��Ĩ�����
������	�$��;��[�T�uT�W N�DU���W{��(t�4�� ��'�t���#��\�h�!I�3�L&)�\��y��х�&�:hл+���į2�wE��>���~����:�|�i��g������CNWЬ�#��Os9�j�2��)T�wa;4��l��vEQ733��'�4o^��6r�D��D�\C�|��(𖕰�����̾�|���u�r�.���Ȼ��Ў����E�S����W{��ܓ1'q���W��uY����v�O��⊲l1�аE��D=1�#�ų�Q�)d�y���n��qY�՚�{]#�I��o�4��o8��3a������t�̢��ƙ��*��g��'�^��4�Z�	�U��?C���T_�z�8\{��"�z�j���[��nf�^�%b�JAi���sn@�9L�du��3[-��?�?%ͺ�o��*E`w؝� �x�>C5�D'&�f�� 4��7�"�	�Q�F$U:�j�l��3��K_�.���x� =����"���(�L�'Fј^�Ò-�b��g]��%���?���5� H8��u��)4,�to�dC�T{u�47s���<���������[���Gw0�9�y�����g���w��3Ӄȸ51g�T�M��A*��B5��3>���<�K5�� +��5?{b�bD"�r��9A�(�R��dLז����Z��@���6<������H^�}s�@��6P�'J�m�^��Ql�n}YZWb=�X���Lf�� �<f�>m����<�
:��;W�XgE\�
���D9��\�W�\*ЖdC�	���g���ۨ�<�(Z�2)f�j������*�H���=A��~0�e���1��)�ʽ���*E�T��v_|Kn���Y9���X��O���� �v�)�xVv2��)�[��%M C��9����%X�[V+A|TR:ەԨƹ.���3g�^�c���D	Х���|�@�n$�v�9��tm��-Wdi�:>�l��� ��4]7X��
�w-bJ�(Ջ�rk��1m�@Y�l���o�����Z����n��E�4���0�A�mߢd%���fQ$}�&|��=Q�6���|�u>�f�]Vc:��.|��%���6��	���m6zhN���ͺ���J%����3S��읞/r�T^�ҫ��L�r
�(�����Tnc�t��cu%1�ٟ�	�9n��k�|l�E��5�j����D�d��TPNG�`���V�Ƭ��1ސG���D���h����N�1HeȪ%#���Y!���Y\�Dw��\�"W��I wrKE�bdm�w���׊L�JG>Yb�4Z}�6 ��|���x���Uj��v�ס�K�«>
��:��!J'����s-����nY{8a�J�8<h�����m�v�Qr��Q��U5�u 3k�)v�T�f0�Kܺ_t<�h���! �g�X\u�2�Mo���l��a�F�]6	�2�-
�(
ȟ��L�%-�0�D�������^�c��*=��+�0�1"�flx�33��?[���))j|��,97; �������a�'����4G��,(��{%.9U�#i�N��Y
{��$/���{��?-;Hn�]��R�2Mm-�԰�)����.؛��?$i=�U"=�#�1Q��K���_=�F�3B���V�d���O�9�<�l/Mͯra�t$.t)�xZ8b���.�@�H����\��d�����{d��S�����,6��Gы�"S�lzi�2n{���_Z����0h*�S�v�#�Ͼ5�p����}��e�7�+tl�;�{b����0���� ���tV�l��������9���u�+��f�mτ�?5ڝ�l۞�����^v1�{=`��Β�~#�_�~Bvr9���kNܜfv��a5���Z�^A�%S��#��e �M���{_�:��џw�.#�Ȯ��P��G�Eu77�(��Y�3M��R{,@�S,���fޒ)@\KuN\v�s����kݥvQ��ż>����Kx��:#�-�N��@A���������J� רP�����2�¾h��ɋ!�'Z"A2~B������/%{�#}�A�;�;dN�1�i���Ц����
qu ���0'
�f"B��H&��k��ӱջ�����S=�I�:���=�7��^���Ć4����+XVd�7 ��}�CUK�)|l@}c���۝@xՔ�i2���0-�W6��w���(�)	p���M�n�oi����l\IG�V<q_���S+맋D#'[�X��*�~:�􊨏��Y'j(�<�.�E��(�L����9A,T���zr���8n�=I�����!\�?��������qSK��֚��������7;���͜�{����~�!hj7$��?��P�k���|�"=����x_�*��y����(l9ם\/DN�=G�-�)Y	��1������18��RG�:��e�|:���	��g;���Wϸ�����71"kO�D���(��EB.S(���d����"��y_��zE��q��k�Tj��7����A_뤝*Is��x�wTp�ѥ��]B/)u�؏�2mv~_��lI�J��E4zmC������ Ia�86_���+&�I��l�� `�N {���R�0�=L���w�t��*�=��C�p;�$V� ���e�d����|�v�L���섣�z�̻n�e�ĩ����������k
����K&?�N�^�l=���Ok1��\��U����(]%2 N�����2�|��������j+!qds�����1�)p�@Ly�[胼���͓�l_�*�~N��_;x���G�*p���=���Ի�,Q���}n��ᵞ��d����ρU|�3�
%Wy� �¾��Z�9��@�Y��'���iPD6a��am� G�jv�9�5Kv0�2jX��+ـi
��:z��ޟx��'S�T�/*�Q�H�K��c͡`��׈�y���N�O���s�cmg�k�#�$�E��ӷPՄ���0)Ӽe�=He�KƲ'v���Hb;�o�T�W2�wF_14V�S�lX5?|o��`��ӵ4��ee��Mw`�C�n<��V��?�Yd,�#à�<4\rco��RW�6$�J72��h�Ah,l�E},0�!�����v+����dUn�P׶��CƝx�������;�����6R{��*۴n�s'�?ƋEtc0�[GK�r��S��H�_2P��|�Z����$D� �\����\YU,���p���c��o"����r`7I��Q������R��V��id-�;9��	��<͉�J���4�� .!!:�H�5گrW���Js�#�6o"n��Fz������R�Zf5�dv# �H9����j����7%g���+����T�K�����:y�Ҳ�g���V��tYr�qPs�
*��&��V�~��ڣQk恌���p⼕��[I��q`�T��	,^��-V5IO��!��;�a��)���$�̢�#��;��XOu\�a���sZQ���hn\1��DȊnr���D���aUX6u�n�F�\ T���	3��7ӛ��J����6��I�A3�G'L�j^*��~��V�?^C��O�2B@8���y�EnTd���4���{�W-�ntuH��a9�m�Y��q[9fz�N�$L��HF2{ڀ�ha���*�݃Y�~�	Е�'�6���KDF��Kl$T�N��Kq��]u�Ʋo'�o뒔Z�[���,����Q�M�V�N*�v�M�TJ�R,��p�{��e-�?MY㻲6K&
$���i�/�b-u�l̯��=�Û0��N�
�%�n�#�6C� ���P��K�+�Az6�-3(����@��R�wV������&yy>�U�ik��;t:Ȟ�кL�}��YƱ�W�lHU[X��V*	1��{ݝ��Pe�ܝ-S^�w�z�D�m-�b{�Ք��uΕ�z�6A��Yr�����Sr���dڳ"�~|��*�D����n��qEX��s���Z�bֻ���S��T�s_KD&���.tw��
]��Z=2q%U;W�r�/ @�މ1b�T�Qijqh.��ad�����iyI��Z�
l��Kd��wU��:��l��k��W��Za%T���eIA)�����t���ww԰Q��6�̜cC7hŮ& T�6-�����#ᬈQ���_m���J=�IRb#����p��䈪.�@U̯����M����1M3' �E�R�밑hk�8�ϊ�B6�\v�m(���߄�1|�?�a��8b��"ŇF` y���t;�V�����|
�h��hN���Ǝ=�d����RW28�x7;���6�AW�����IJ��e�()�ӸL�L�~�"H�_���I@h�ċDRl̮m��lM����{�e��:���U@ͩ�������.�b���t�X�h\���`2a�zmY�A\_��͔>��G����f��{1o�zʜ#$�oO�Uʾ�  �dA�X|k0�D6"BEDZ�_�-�ux�?��F��:^����m3��8ӵ���_��U���Dx?	�i�+�,�����4�$�#�
�Z?���Ď�-.�������P-[ :��utn�~�Rb����Hʖ �:b�hk_1��c̶����
>�G��{��Qe��%i�Q�^1ھS3YSnH����66�@��byᆈ��.��e�G��	*��#o�٨���#��9 ɿ���p�Ԫ���ǹ�.:�d�e6>�g_��l��էvG�R���, �#V��\��QG��Qb#�1���Vz�6��p|ȻYK�4����fN�Iȩ��G]^/���^(��)*�v�Tި��!,v�+�`p�l���k�Œ�K�j`81j=ڙW忉�m,g�&}�ɟ������m
0VͽÅj�NRp�Цл�%_h]l���P�h��.{�_�t��u�ލ�|79af`�#'?_m���pan�P��X�u��'��h]MKG�3�mVD���������-�#uw��Os�R�W1|�o�7�k��y��ϒaE�i���J�A�d���Мs�BXW���.L�xO���l&�8x��V��}��d*j$ȋ��ۮn'���3k������QgNu�}��1G≐�XK�����{��ޑgv�Vʹ�n�W����%n���d�v�ij5�{��NѝU{9$-\��������-���[b�	9K�`�u� {��EO���w)a�)���\���k�6/��K���0�����L-׼���?���"�M���ZpR�e����٥��rd��Y�
^�.@�.�̻Ә�N/W���Ou/�X� �gv�0���%�_Tr �EC��!���fU��u��`���"��
`�މDݼ���e��SG0+������qZ��,������I� ����[�
��-e�]�oh��nI��憥 ��ىP����|�0�8h�Ri=Ew�X7*��d.���,d�Ηz�+r;c}�@t�������F'��4㉑ޥ��ѩ��E�K8��-l�e�J���@�bu2tn�bv�AG ��"et��R$T���K��GP�b�\i~�͙��6��� ʞ~��c���馦��^��C�s�N�������M����/@h�!pG�1m����0�O�4G_�I�@ ���7뫏�a7��?�#��Mԍ���l��Re{N�p��>l� R�χ��KC5S��
6�x_>�O�c%���R���d�:4��������R�cӕ�5z���1��f]Z�U�8�zM�ź�Pfa�̮^ʱn��l����j{S��DuϨ����f�.���e�+��Y&��:����t
� f�1�V��㹄D0m���2f�U��njD������R]]DX�ڞ:5�Hx,�#F№���E75H��	���'a�n�(���y:��5f 7��m��
	Ò��!b��D����Wa�͢��zf+��{7�S���>-���>Wv�C��43�[�wc��H-0\�xER8�1	���"������+�2������W�%�U��Z��8�@�w�& VHko��h�)��;��|+��f���;��u]��ߩ:���ȭ��s%X&��a�P?��R)qw�ާXb�A�<s�a|����Ǝ�,sB�����;�'/��H\���̄C\j�;�]p���:ǎL��2΃&�8���g����Ҏ���i3����:��p%'�����v�a$�H݁�27���J�?�GP�X-���k���?�!���NVu�d�C[�ʬ���UG��/t�l��3�M$l���<_|0�s�u�~�e�gy��]ʅ�śB���у�c��d�N��T�p�ۗ��>!]�uNm��$M=�XIzݝ�K}b����el�ًX�\�tAV䆝i�AA�E.��<��
H&�hY�*��V}�<l���م���KZ�uV�V*�����ʴ�{+Hu��c���N����=@T��F︶}������W����G�)\�Z�=rj�R�/���3��Y�64TO�V-:|�u�����Xո���_e�f@�Q��P8/?׬4R�Q���������9�D{�$U��х�m~̵�u\J�Q;=y����%�I�Zm1�1R(g�թ�B%ŕ­����(�P\���@�M��ە��1A�
1W/����)��~���B�x0�C����?�Z��@ao`S�-�tj��,�	 $ �~t� ;�&��{]F5���q���Q������|_�w��{3�,�hq`�.G�;|�F=��4�^�vve���l��G��&�}gȷ���kc%SV%��:P���&3g�շ��R�`��4p�9t�y�+������q+�UoODf<I�`㖿g�`:3��@�F*��6
��k�&�6��б$���-���-����}�sgЌ]3�������λ�#�@�.����:��n
h�	ҡ��7��X�oK����4㫶qUx�T�Aǿ�P��Ow0ۮ9�D������{F�ǣ�	� _�]�rZ�U���0�V����?�uj�����&!��!|e��$�x�<?^$�Lp��l��,K�%h���=8�ec���5�끈:�i�0x��!�qV���K>	�4����j*�-ۙ7
rE��hUʮ�����������&�IU������.]��A��˶���#)��0�i#Σ�	�����F���e��
0ux�XH[�*�Q��?$l0п�(�˜�g`��j�C�)H��d>-J8N�����2������ђ��>���7j��X�W�dI*e\Is�_��ŝe����)-��4��`�� �0 �G_85�P�Ƭ#c�;��/g��Я;4b�7f�ĒԼGP���6+YK0O��=��f�Z(�x��=��3��Y��+H�K2Gc�} �jU{��r��K&��Ȅ��G�SŝS9a�Ɍ���}�f�p�)Y��>�i��_<_���!��0��l�<2�������+���X(�}��i�?tp����B5MQ�%K�s��(5�	�Ⱦ�Ew�t��夕�FZ;��=(��C���5�>(b3b�J�����Z�~+�%�+�.s�@a�!��>v�׮|�~A4�}�,Z�D�8���_�����42a-����&vwyDk�[���`�8}� �>�4"���k���^��W}h�|�/�X��0��K�8\�@��B��Y�F�����k)ك�$��e�~�ӟ./���ko�3*�'�.�D��}1�'����7A�	]���[u�C(�Ds)�PwǍXJ1�o�'|E17�Բ�ۥ�d�j~���bM�:Xd2�&RP�wa��Q*�H��X<D�zA�o
>e!^��pA�.qY}����Y}1J�l�I �d����ŷ0�n�?��}��$�J3����~t�4}_�O��0K�2rj��لNp��}��w������qK����xR�,'������]y*�bk@���R��^�َ́9��P�Ōv��g!Q"�d�mn[!�6~0n��i��O4�R�����{��	 �h�&�V���\mXQa["�����RN8;P7gxŊf���T��q�G�V��re\���K0Q��ZPP;0��c��66-x�-�oc�&G�|�����~��Mv�2Y �t_V�s*d����#��侃<݄v�h�Y:�
:�?���`o��"���6=���m;�����[ŝƲ�g�C9.�\�$�:JQ'r@c�"x8��ըo���
ɂ%����|�m�-B�����Ϛe��<��18�<���HiF&�w�V ��\|0.G�/:}坿��<ԇ��]�ZK@����ڛ엢��v��p��}��ޭ��<F�뾞�c7��@�|��IOl��>H�M@i0^2�^ǻ�� ���J��T���D�st��� �yI܃��I���8�c�nP�ַ$Ce5�^�(t����{���}�^�T[W��Z``�:/p�b���X6����q��x�x}z0$JO;�9�kT�27�͙�C>)�=P��y�=���Xe6[�r��o�O���	��!����;�v�Zh�YWG{�s=M�F��>�E�n��m]f5=yVĨ@�c�2D�f
u�)����^��JRr?�.۪�dq�~����$.U?6�;�&Gɦ��������0�a;5�raׁ��iI1����L&S���P:1��.I�Tm־�8�o(��T3 +^c�NI�kyi�
��z,�e�d���x���c��h����D-�o#H\�7|��bi�="�בX��^m��R�o��I�]a���s�g^ew���!�R�/Պ��e���SYpȞ�����4�Cf�H&��'ّ]@�E��S$s�VfA_`{���頠��; �K��N�,��v���,����/�dq�J`��ҕ�K�o����M�n����k���
���� �L~��i�T�%U��<�t��v>-ͥ��=e��Zs��N�jKj��u�[r#֘���U�d����V�i�y�xk���Wওp^���Ɍ���&G�������$9 �w���t�*��ɫ��?�d�!��	��p���A��lvo+r��-s3����JThh�-P8Vtэ�ՠN �(m��:��҄������3�u������;���-wKތ���U�U�=$M �a��HC�b��fui>���\�������pxV�C� ������F�f�(�f��U2�T�+v1vf��b��-��m���Ru_�1��5��@��4�
,|�	t�KD>��gC�:`P�O�d��T'��@0�����>Bi~�m,�L���������8��{X�����g�⹷��^��
�!o(er�o�՝��h�S��cڿe2��q��cX��g���d�n9*1� ��8�ɐ�S(���'k.�h�(9N>�Aj���љ��@��?�`�~m�`��K]��;�ةR��@pٝ��p���h���k�İ9���D�`M'�0pY��[b��1����Q¿�߅fy��Az-_�#����$pmɒ;�66�]K��_��U=��D���a4�gC�������p�'����U��@�21�zS[��j/���Qy�d?�_
I0��,k�ތ�QO.WXY�`H�)5��3��~�\e*D��,i
�\Q�bNd������-�������F��w���|���lՙ�uSy�Yci/�Î��X�n��u+�a�kq����?_�/��(�����"�	b�~Q�ͨi�g#s�$�=���Z����۔��AƤ;s:��T$#�{Q�TE��<u8m�Gt�4\���$��ö0&���m�m�H�3�`�>�l)c���s�0PrC��Po#��ӬX!���8�v5o�`RH��]���꿮����N�������I��~�+`	��r3��0��^�8�S�����V���4v���^}��&x�O�z���"�r7צD>3�@d�"�&9�/p�X���d�Y+Xj��f��	[f�{����IM��U$&��7Y.6�kt����T�3̧S���&6�2d�M�ЊoDTN��_��(Ζ.{�����4�G)I�sI���F�����2'�3.�|W�~D����u'��ؖ�B"ZdM�H�+��Ò m3ś� �gu���D�"���$eKw�����6B"��Icn:�d:~K/	�с�g�P�JBl,n�Z���縈|�rNc��mw9�����O���S_�zN�����O�6��C��7�3]�ʥ�J�#>���j[�U9�j�s����[�Y�M���*�(�%������e�"!�O0�l��F����)(�wM����6`����P��V��0�q�+�]�xh�&yD����`������_QgS֤Vӡu(W��7"_�by|}�ވ>N�G��O<OD>YOO�z֣��*i�����#�	�*�0�8�@2t�7;S���/��#�
�4�>�Pm�v|�J��E��@�FL:���z`�t��PF@B�@C�[#(�?J��!zqo�M@(�1��=���롯�g��Jyw����MqZm�"Em̨�~I���ы!��6h�_��Q�R	��H1)-K�eB�^�fA��
�%�2vY�u"�oO��%�ɨ�5u��DLگ���~eqE���PMx�%��寺����j2z�sd:���� ts��W���9��U�d�t���x0q��"��g���E*l��/�������e�T��2Mts-]��%��2�	�s����L.$�2|��IBo�]��-��&��˜��gI\�rPڅ�Jl��9^k�L����Z�q��%iW�W�rɜ�-'�%�Մ]�u���jb��֞�8�:�M������o7zF�9g0�9W$�-��́���Zi;l�B^��T��������/�ż$*s��Ii7�ִ9�ț�K����㳙0����ΐ�L�gǴ�0������+Q�Zn!�?��4ʳ�V�T^4��$�3���9셆�l�~�E+���CVC�>��s �f~��e�֋��� �K��XAQ�J�hŜ������\^7�nr�ײzp43l׾��?��\~+����ΏoސbY����|e��ɬ�Cp�'���Q�k*E��d\��H,1�� ��+~��}�p�0r�)3S�7]���^���
�st��Ua1�ZNQ�C����T�O� �s���8�8����C��1T9�yw�@� <Z�����]�A�f���s�'0	x ϛn:��qRLy3��e��G�q����t>a�[ɫ$;��}: X�ȸ�S�+YhBdx8i�S.���W��`�J	�G`��y��0��;a,�)�Q	�����$+.܍��0�J��fa�/�g���Y�@|���H)i��H|�B%�]ۛ���큜f�ŷ�-��J�"ǎ�)4�\���}[�;��Rh�,9�)�"�3���X�p��=nf)�N�yK�E��㌟8vU1V+Z�1��� �������`�B�'��>��7~����)9�ʬ���d��hx�k�:�A��vci7�!4����/<l��Z�?$v����Q���+U�
��xb�k	�=,;ݡ՝�FL7}�H��P��ۃ"k�5r��瀨y�=`�c���V���Q��ϥ��_��q�n5!cMS��］ǉ�ݶ,;�P����n��r.�ijh��,�v�cJ���%+��?�8�¯fL�"�\���Wf�s1Q=Y��}��w#����i�8ya�Άܿ���Dp���Q7��G�9|� �O�W�xY��QdE�����Kx�a}{r�o�<M��R��L� ��2��o�A7�%�=��P� U�\Q<]��aO�GK�+MŪߜG�DT��3g�F7)��20!C<$(���i���N��&�w7�KH@�m�}�S��+�#�}���1�Y8㋷C���>f����-1l3kJ����g�g#���# �����9��f�z��xҏe0�=�eS��R�!$/�Λ�QnI�G}e���u���gI�#�d���Y�8��WɊ�.;��ՠ��y�����O��X!o2���9��N2�dkf��C���7��*M
��_k�	u�v>
Mǅ��5�������K��5�U��&������pi��5x^6%�(�|���	�Y�B�[wڟ���ֆ��4i�PC&D,]8.�P(9[�w����eLա�N��UIڸf��H�f��)�唸\%�tECh��Y§�DX ��K�ߡ10��@.k�<i�U����(�a�jV��8ON +Ͱ%��oВF�=~�S��C����Clb��J�bz�9���`]+e���E�}�k-�+�9w�өIU�PHd
���i��`j ���)r����mg�̦c�y2���}VPM޸�k,��W���bv}�Avb���9��w��k��t&�4����4��7S Ϣ��C	4F������q=,6p����|��N�0N��"���t���&�Tq���l��T.�Z6���d<�"��i��VB�U��?� ��#��d���HSw���4 �n%՟j�C��%��
yGCE�K��[��ٷX8��͵�/��� $�EsZ� �x}��F�K�J6*e>��q���q"��3��@I"��#k*��2)˼m6wVE�PDp`RP���f粷�k���Z�|�
cHJ:5��?�zt
��]a
����`p��Α7�����W�4gD��<�n/V�����E/���\�	DB<@��i�Y���t;�C�%%��S����R�x��:*�Agh��DXE�o���/�~���?pm����^��%g�V
v&׾$o��Tw%�$��Hp��Odr}a��^���A�-���1��ʔ�n��Eb��]��&�Eo�o�
.�"���]Pł>��*]��hl_%�R&\/p쀻�#N��Qi3���zZ��U���bN��?�|��^kg����8�GU��荆IS�WG��H2�`�J�I��|������m���1�s�����H����o�������z��(�'ک�=�+�/�|���2�X�[6}O��N1)��	��id��g�7ٷ���{A�@AAfg��O� ���mŶ���H%����:�O8?�`'��xi�Z{F%�N`U��O��B���V�]��C4��Cs0��0��%C��Xt�y (�1��l� y*u���|[�ʑdCέ��8	���z�V[�	FZ*#���M`��ŚmЦ�S"	���W�nsܵ���e��~�et����Q�+?��-�#j{��.�fz��(�͙G��I��^UHxM}��Ƈ_QV$�g�� �z0E<]j��qe��a���q�:���~0H7d[M�1�jI���E5,�)�C��¹�>���z�D��l���ٽm�e;R���n\��8�S/��+SAu�b-g�)ɳ� .ʙ�K���ex:�a�g�0�;�brd���k�	���� �v��s�	�T���Q7���~2�6P�~�������#{����y\I����|���������+M�a��Qۡ��<�$�yM�E9��}7��LECy��x�i���)෮��E��"v��5�[�*�&'*�<YB�3���ąguy��>���0�B;_L�	ƌC��:�GLZ�[���5����]�`��^M�.3��ʻ���˅�����T_({0B���7_	��7�[v�N&do��.���PiG ��iF����m�̋�������Z�HU�zz+��['�V=;$�$�s��;5�;��VJʡZ��@G��}��a�3�]�_:�cE�G������2��h`u�}Ub4���ˌgH��� ��|9��3@ڶj9�\�kF%J�'��P�2�i��T�l�neW>����o�kTȶ��v�ߴz�[�����x���5{�ai|;-BX��ʺ��4�D�������$��mFn=��T����qTה:=��+!�:9a���h$ݭ
��S�t������!{�����qp,[��@�#����0�W��J����06;����E�ې��i�	�M㠈�mhRt�,=�ޑ;�Q�Y�����ki����u�A_�Vخ�q�C���g��3�P0a��l�ݴ�9).�icn��ub�L�|7��ԉ/TZ�i��-��w���>�ĥ��;`Q������p�Ct
n�g�P{�Z5Ux��WYU�BB���<l<h�î�!	4�=�tuq~q�� �v�p��L֕�vU�,Oj
���;�8�u����,T��,: ��	<^)���x��q��D7 bA4��S=���q?gJ'lEd�F�_���h�����Ur�󹵧C�]扄Q0�/-�� �N�0�x�җ�	��i!���M��'�J�����p�M��J���#k�n~�����@yZ������O��vv���.2�.JY�_�!,�\R�G���9"��nyS4;��U�	�#T^�=�\��jMw�m�4��̈́�C�zcF[��V�x��g�9���'��t�O���_E����s�ש�7�VmR�A�����!��Y�ı�.U��m�È��]�Sgn�L�l�#�#*��Q;��},��=ଟ�W�B���Z��&
C#;�.�1{��m���9����`�&��f���ޥ�B�߯�����ݧ\Q���q(�m%��u%��`�� JY�.Y�2������~&N��ʲ��<��>EpQ�Z��|�'����}ا�_U+O�+���o9y���֨×!��@n����*���w9P脹#_��b iPK9��|�Κ��[T�s��C�|��D���(2C�
3�$Und��3w�k�D!]ѕG�5-��I]���DV���d��j�'2���we����mh�a� �+��<��mQ�48�%bym��9���Q�D�*h�?q_ك;�B�Qo<5��&�S�un�'�#�0��W�����e�v�y䊍�tms�";�T$b��G��9���#����at�uU�~��6��-?���L.�Q��VH�a��H�����f_���_���I���.BA.V��+.��걾a�&K3�� }OU���ߥ��q�OWJ�nX_Ժ�/{�~FPy��*nE�fwu�z׼����:X��Co�u�Ae�]O��T=�uNسv�$]�N��i�욼1�qxi�������!�Ǎ7/�b� ��4�����P9}�B�/�^�g6����b�Џ�!Z�v� R��i9���3�4Y���P�I�:��!O��	v7ׯ� NHf_6{9#
"e�ߨ��#��ʪ�����r�O�p^ -)�,��	�r�2��ҌV؉�A0�1a�|�Ɯ�[�/n�m�x��R>�J�N���|���m�@���GG5�Jg��#eo �J��R�:��5��g���o\|������!�@�9�%b ��e{���^��q\d��YZ4�xwז_��0G���1&��dʖ L�E�K��V7�P�r�]��
YkÄ�H�!Cg�؎A���
�]���Yf2�xVZ��?��2�{j/�bZ�cơ�
�EUJ��gv'�P������_��0�&z��p�2�v���4��*�7w�y{�$���N�1���j�W4��ɷ�������^�2�5���?�n�YK��u{I`��S�IL���<n��n�T|���<��	H"�f�'c��ox"e�X9�x]�.�*߷��/�s�;u�m�y�@�E銕b�Q����@��&���\�Y_��"�vIb�7�r!? ��E�i ��U�u;"�/\7̈́�Y�_z�t֊�
�(�����s���X���s��������hm�#�}O7����vF~Ӷ+��&e�[�l�Bm�Z!�a)����L^��|qQ�b��Z�MP�a��R�2��cDM��%n{O�����n�ڻ��T��+�}y���g���C�}3e'|j�u��5ꈽ��t��)O�F��{�J$F�3N��,���n�i�_�g�V!D�(���n@R˿�1�;c�0,\E�2�cZ9�[CL��%a�P��j��6��]N�7�R�ĸ�m�Wq���L�?O�|�%�ޟ����WJ�1 c̙V�����Z��b᯹�>��6���4�ߓXtLV_����R5�Ə(�/~:�Y��qi�/���Z�:�����÷>�*��i�"F�ɷ�暳i"&wKLB�������@�^���%S�?��^Oۺ��"
ԅ���Z�X�f�1�Q�x̃m��g���%5�~�)���5�4��>�Bm�x�?0>�E>6\��:�)~��o��G��6�"����Ù ��7��5�� �p�p)8jЙ�w�N���8�*Pɏ؃l���/�� ��U����h"�v����p��̯�2wyl#��*�-`X�&�����*.]O�����{��2��F�x�'M���� �LUn��}�>T���H8.���STZ�*���Zˇ���"��z1��ι�s�:h�G�/�}-�{د����[�!�� ���1U���2�Z�Eqsѹ���gwކ�(�o][���$�t7��nc�ӡ�Z��w9^�*|���4�V�������p`5�m�tu�`�wMX��`&��Ji�t��m�� ���,��F��2 ����}�NAu��5��[�`t���ُc�����~���D��|�se�O#"j�N��Z�3S~q�+Hɑ���Op�_oH9����I��*�jm���tQ&_D{uDb���@�8r�&rQ���v��Bc��:�U�֊�3%v>Wn�rS�k
���)� R�tU�AZ$��
$<:�[��M�˷�� |H���ɏ�L
��x7�*�r�4�=�1r�E���Z �/�R������ �F���-�Į�=W~�Sl� ��Kq\	d8{��XEU2��c����)��4M���-��!����g�y9E��?�k� 4� r&�-�m&�u���Gڎ�ں ���c�́��8�����L��� �M�T0�Q�O���h�^�U���6�>���s<��z� ;�cF"Э�3a�݈z$��x��@sj=(Kn��vޛ:���w��k�o�S�8�jAP�[��;L�Z2 �7�O���� ��)(�yX� �t��̏^�|%���q�p.(v�
�IrW�����K��y9�W�-R�����̥km3��#TV�2��B�lщ��.M�}�h B�T������H��%S����A��kɿ�F�>n�W� ���e*{�d�cqMb�4��>�Kܒ�*+�`k|����g����:U��Q	�b�:k�0��gի�äB��V Y��R�A��848g�%ܓ	�m��̭�Ɍt��ך:2!���f�����pC~�"�*Б�EyۓQ�ٟ���ͭ���Q���N+
O˾�ƾ��7N�Zk��>=����\��v/ ����RM���i�����PU��9Z�f������y��h��Ӎ�Z#QG�:]=rGz&���6{�\��|Uh��+o�t�_�Z� ������G��Y�PKPH�7?O�������ɥ�4���Z���e��K�;�sZ�	\��Jywk�;�/mi3јdii�����+�0^^�����~�%�-�0Y���ַ�5!M������WDݑ�N\4������g���#�2�Is�iyru.d�s�Q�=�I���kB����z%���<)Uy39Z���e�������ɣ�罳g^p�z`�\Akm��{���_`n��0�`P6�T���k?�<7,߈����1�hh�F����ݷ�zMUJq@�V6�7:��)��\n�d��;j�Nt^���3�"vY���0�9�Y���ݾ%��b��5�%'�@< ��iF��tӝ�h�k��0��,��SPkY��d�f�K�4��F\!�/�drrBt:M��t =���1ګW��W>��C��rJ�֭\,�Z����w�[�����S�U�p��]��58�iX���;٢���}n���3��?�.����P#ԟ��"ܲ{:k��D.
����A��޷K{�w >�b��6O�!9z@z�Ø������ G�7s�lʉُ�ta���-�!��җ��#�?���O����	nB�K�wOG��Y:�Y�V"�'�s��ZĘ�{�Y��g��w�%�P��o����0L�����N��gk������v&�o��zn������S��U��q�{~B�y]W��s�j�X�>��4{�	I�_V{�^�Ѱ%�p�,�`(�����T�m9E�Uj��Y��ۣ��њ�
���yD�m�����8+��pU�q����;��@�Ҥu����gAC�<;gI�7f%�me�;K�(�i�>��v�.�|Q�/���Y��]����n�D��P��w�n����ʚ[��E>a�e�t��#r�6No�E�)��X�C�;���������vf��7%|��,W�_��;8#����kQGYe��pq-ۋS���?�2Q�4�4��}�}��|K�Y��d��
hM<��*���u2�Êz��K���hV�����!a�a��Bj�,����X��=2ŔFU�S����S�kZ��ɕ������jȠC�K�$}�I�G��;"�OedQė�u��UV�]�Xz���Ba����8��qQE�c��ܽ�u:B��)ge�����/���x�g|���G��o�FF�6-7�8�jP+�ˋ�J��lX��BkϵG%y!�#�O���������HJ�����~��׶�	 �{�xʐ�+�:J��*����Qc��w��Z�J��E2�"�c4-���_*7�][N�;K)�U,�\_s[0����z�I�pQ߶L9>{C��k	Ŕ=XD^�qP/Z�|��bm� #la�a������0��	������G�:�	'��%f5l�=� ��W�U����Nk���XC���opG�x��>'�?�k�"W���<k�O����l��q�%{���<u��<��CmU�V�Z�{k��Ή/�W4�̚M�d_o�s�g�v����J�L����VHLfS�g�@����V��P;���O�������f2op"����7U������R�mhZ���;�*h��n��#5�I̳(W�h/#Lx�ď�$�Å�'ݵe�����;ހ�w[��� ��`I_Xކ��`f�+�{���C�-S($x&�������w�	!��4����gm A��k�(���B�*�u���@BK�[,�L`�뻀�Sw6&YU	qZʵa%#VL+}9HINl�D�aή܎�d�.�	0;Um���ý���������x8+����܌U���ѹ�DfPk4d���6�%���4%��o=s��YΊ�lG������0M���e��W��d�z<�3���4˱jg�d�A�:��9����2ES	��d���8g1y{��XU~[O��)CGJD)i|de0�J2�`��<���<�@j��;��IՕ�Р�@"���N������'����B���^(I ���H��@< pd��ݾ*���4k*���
�ܾ� �g�4EQXto�Rw/.�R�8L<�Ҷ&S��Ċs���r�kF����җu�alH�:P�b7j?�j2��~(5��:V��-r���`����q:'���GTp�@-���+T��(����wQ�î�^;�B��b�K���~2��V��P��T�0n|�7W�6�P��Q?�,��ʬo���k��jWH;�Q�(�h4�̾�R��GH}�m��ﭤG���u����t�*6�Fl�)7��S��ң�tMi����5�� �]@�3��F����� �2��m[ˌ�e�g�T&�4��	����� ��LD�|*�dYn�Ä��;;�z�{XM�Ԏe˄X����ߎ�.qANl2�YWx���Zt�%\��qW�Aґ�#��!�t��=�+EY�����d����3���bQ�?�ܵ\�Q�VL/�h���Fܲ�ד?;�4�e��q��Z�O�Ȓ�'������:�z��c��D�+�"��Q(|������!&�N��?���~]Frav��`��Q����g��-}�s�bX��G�����S��W�y.S��ְϝ���:`�'LXEKb�[>��-����0��2U����(�Q���S9"���g���_>��(����IY/���o�M���QT\ἔ��O�qZ�#����`}��*~���A�'r���d*W��ѯ0�Y��Cɞ)/-A�̩��A��N�^����!�6����f%��{V��z��,P��v�X�È�6��O�Y'z�D��?��x-б�����H�ۮ!��fu��{ 虑�
*U�of~0��� �$W��	@��NG1=woݏ��﷑�������X����A0e�1��&�}�r�F=
Q�� &+= �{9��T��M�kB������"�E�	:����k�%QX��s�%�/���8
��>�~L`�Ra��[�;ߥ��KP�F0�jke�?|��,R�3��R���5IGfs(���=Wn��m9G� Ϙ� a��5��>h��!c��,��$����pD���^�0����5#˧�p.�u��R����XGN��J���3�]z�[q1�i
���hk�f7Kn��eV��O(z�#s5�J��f>����wo��la���@�g({n�
r�E"����3Z�q�6��Q��KŢ4�a�B��<�G��h���6����e/�YP��LA�:�P�б�Q�kB=쀜!�&���m��%ZlI��¾>h�#st c\^c,�p���4Uؼ{��f�s
��3<��_�Om��B��G��%Fa݅V�"�"�>�[<e�X� f�,��3+���肻�]r���2Hz�#p�͸�:F.r�]Cʎ����=<�;�g�'�z��C�������#���A�3��Ho��y7�v"6]���3tE�GX�^�����[����ƅ�_���#�m���
~o�9�w�'}�F��f*9�c�$��階36�	��0<O�+ʂ�!�(R����r`]�����_K@�
t!,eZǒ
q�KA���ݓj�Ι�A{��8�A,�G|�$e/z������M�0����H�CJ]�`��,�˕-kq���`ȖOF�g��>�_��_��K�#���I�{�ٻ��zL�gYfB�cD�b���j�N܅��?�FHf�͵zF�b������ntkы��e.���!t�jaۋG��l�����^aW�z��Ze�u�ٙ$s^�)g�;b*f�d��9�3�"ܘ�gV�;Ia��@T��հ��ҙ��k^n|���:l�UP�;Sx�웲��oݙ�$�9�=x5�|�Os�;���u�����g9���RU���5���I%&N8���aBp�Vʳ[$9T\��q������x���T�O��~��˜��t�'����Ve�Z������$��A=錭x�x�\���.M��GS���cWS��	͏|��?35^���u� *�.ؾ�>�����ySC��A(�F��|O~�[u0�IC�g����O�)�x�a*���'tR0��X��������8	�b��b��ZX��gD$�V�!��>	�H��i��,5�MfjU'��1����[��=�*�}���t��0�[c��#N*b�_�^)��(�8&ᘚ�g��h_$����W�jt]nEtR6�Uq�u$�Q �T�tf�q�N��2�F��1lA/��Y��m'�_��<c���&��&q ��lg��I�n�a�U�]$�wfD���qzH��=��"��kx���O��i�������T*��
��M�w,^sr3O.�&���.���!G�{�]*Q�O��\���b�]��ڸ�+��Dh�Q���Q�!��V�*g����I�UQ`��G���%E��n-�u���Ρ�N9�n��Źl�6ecn'F��LCx���~bP��Ν�N33èΜ]D�K�90D� ͂�7ꅕ�(�0��oA���8��{���_M]Y֘T��%�h�QO�c����7��s�nbRY{2����p҉��
�J=�IM�1^,"?�P_�N�>�����5Ġ3�j��}&l66�ΗoYʠ��{O�ԓ��>�͝.i �
3|��fW�]�(��[V�#���UOf�g�W���[v�x�!
h���U%X 	�JΞ1�w,e���s���Z�T6G���$_S�9�D��kV��R0�\	W���9l!_�,6"{��5�a@wm���,�׏�(���Y�!���Dxalx잶��z�K����2��%�J�M5K.F��=�I�`�{��3��QY'���h΃�� +�ޚ��E�y�[��+�.���8ɛ�8p���C���#N�m����y�DO��x�A� J�`���F�!d�6�R8�8X�_�-��tMfh�h�g[3X�An�;Լ��L+!]2��]��(pg�mK��a ��䭨W�I�x�àD��O�+��+t:
��n���`���E�üXi���u;�{��Q���"�2���'���ɩ �á��g�d,{艟Yk��ZAU���h1[q-���(
�Y�흥@dFnPRS����;�n{�@ܑW5VC��,!�BCع��a��ĥ�BS��Q���^�E)�d�S
�ǽ�8��C$��mlD?��с� h������H���@
k����ѓlM��>�$-�s��T�`�f|��X��[�rKDǔ�	E�u�{��&A� y�ݧ������:*?/ۆ �4T(��tj�Qu�A��!a ;+j>,��a��?�iOp�Y�;�.a��b�C?8��[ ��v�u>��ъ��R�h�[����h}��R���Ɣ������ڇ|&"�g��3�J7PC�C��PCT���SL+{�
�5�@���7�4�{����mC��V��1���j��A2֩��`w�-h��֠��g/A^Y�D��|[D��i�-z��uc�;�\,�ٜTSy���x}��;������e$�������'������Ve��;m��#g���d9�se��o#u;r?���P���d�4�+�i�����f��u���?C�	�N8N���0�;)��f���"x@$W���s��W��%d���!V��a+]jڑ�5~���tm��7i"�O^l�$�����3x�����o��ԁ��=DI�_ �N��)�$�j�3D�2��;12r?\}擽|����m�k�SY)���{'{at@V�F@Pϟ&5�IL�3����Ńj��2����:�g�)E�����m��E�̧Hē��:���K䇬������fD�3n��=Bpz�eE]�+-@ ,�?#]�i�a���F�>G�D Ѯ��W���6o���p�}M���M��(yH�ĠB��`�?WID�T��D��ڡ��Ⱦ"�����c���`8�[G�f�d�����sJ�&N��$ �?!�7�}B�
��yn�E�h4�_;X�Cz�%&Cw�0m��1�����!�����Bv���#�ccP_�72r���m��L��*����/�{�� -SGߕa���Q笨v��_  h���Л�����L4l�ĭ�T���!%�彭��L�i���P�����d�S�q'�e"�u܍�۳�����H�B3�P%4�˪t=G؎�d��X,%��'�!��Q���`3Fs~�m�/����S~/�TX�I�k�N�
�%�d�fnR�R�9�Y�[�J���ܩz}t�&&��w�ԀM��OI��>_�aLeYUDsv���Do�.�-��\�L�U6�$��b�U���3�QA���!��+�~x�
ZH����@���O�W�Aj�5@���?l�	�$��8��k<`�}:p�f���kʖ5�V��q?��×��9��b�B�!��T�
|�I����z�km>��;�u�0��������(��������v��G�T� ��;�ȓ7/8NZ���)��o8��{b�o������9��z�רQ�<�$a�;d�U2ፆ�3��zn#;�K��J�ocL���W<o��"]\��������Jd.r� a�K�j,��� i:��w4����#n�r9�숇���*��Ŵ��*۔w���!$*de[#H�J J����V�x�� �:�RW*�n^%c���<��V�덈`dl�1 qt5z���U����	�_y�[X^�۔���?-����=
�'�U sfG�������`��QQ_I3�j�,�8Մ.����<=��0NZ��&ݫg16qb��6�/4�=��b�7y�����ɫ$u^��=��W�ȿJV��$p��/}bM:R�!��V�lv���/(�tx�z&,T�W���@����P��O������P7?�<����a���W�u�;D�Y�]��,�����W �0����ܗ�����ADq1z�Eq瀑�s5�;�F`����?��S��`��u�aq|���:�M������zx�xw��},�`�F�2,Lr@�����+
Ց��Ǥ�z(����ɮ"��8������5�B���"̋��#�f�U/|R&�lC,/	8l���m�P]�C���.2}B�������:��`8&D��c��f���F�jg=���M�:=%��(L�!�zi����_M7�@�l3���6~�s>��Q2�χ�33\k�h�V0$�_Ϗ/�,�(��S��b�U� LF!������l���� ������Rm3�H��'�[daD�][�&q��p�K+�!' r�k��8�\2�k��.9AX�8K���е��`�����0�Ѕ��������(m��<� h<����#�A�3�L��ɏ	ɴ.�kR�%Y�>��纃v刴�f#'���@�(U=Nw��5;2]�Be��x���b��s&���HO`�E�8d��1�9u%�"^��.����s`��f_���	ۉ���fm�m�cJ; ��`ňRB�ZP�˄�f+��C�^xA�$�ni��'�5����}T#C�G����&��|v����4�J�CE��^�v�'>=���?��")���TX���VAB���ess&�%:����'/V�f�m��)lf��s����\�+��s�$�b\�*�N SA� ��AZ�ٽvŐ��|g�	�y�T��(���y[�P(4�(���xN�7!7�xhS�EoN��'���_���_��.����r�n��K^�|i ?ڼ؎���9G�6^���:O��0/;�scZ�{a-T���v��U��񒩧����|9F��䘘��G� w��q�mJ�Þt���z�p�q�b1' �g���.�Vw�5��9d�s�jH���T�Hjmb�I��rk,a�<���؁G��:�;��+��;�N \��E��\+��0c?¼��Xe+�?2� ��}N�bR���{�nf_)�_��_��{�J������������V"�U9�O�h_&�ˆ� ��s�4C� �&e5]#s6$��y�y�ϓ��9<�z-��~�V��Lm60q\��L3�����|�]N��E7�>�_�74�2V�na�����҇3���iܾ���=h!��<f�y�I-{x�������" [N��)���Q��<�+���	�,���|S�q?u��
RmFӻQ�D^,Nj��v ��&�)�.�-W�oS��
F�FЂ\��ȆCW�Շ
�^�����kh�v�Bq #��N�k�#���w8d�2=���r'�P1B�c\����+������d�9H1Um���TSIyh~L:��c�K&���m� S�nZ���d[j���e�*�)#l�Ld����t*uda\:�Ɂ�F'w��T%Sa���iY�}/��I��k�ߥ����`���~��h�k�,�,��Yy����3��k�4yT	 ��T0����l"1��&"-��`��y�"c����kR�|"yz6A(Gv?|���J�S���3�:�A��_m�9,�����[��VS���Ea�<+�#֫|r(@��"���]4Pxᤒ��nM\��$
�Ez�-���N>f���2���.�qE��dd�6��E����c�Z��R֫��݊�_O`��K��*����#{]{i�AP���/u�Ŀ�%��U��v^�
l�p�3�>x�ӃL+�q���~I�熐�c]"��
c��=V�F�I��k�������i[��=��84x3���ϐ�7'����
^�]]���~��7v��A��T�G,t>:X�=��&�]����Ma�>���E�\+�����M��ӻ(�\u�j���V<�����^�e�*d,�ؘ���-,�������� �޼���'�����P6�ߒ�$��Q��Rf�@�0��}�d�u:���<�����d�XSh���3Qb77�����z"�ɭV0,sr0}�1Rt��'�1�t�Q]���:�[�X0�es
���r������Ne�����v��`���	�\G{�N{A:\��=�Rv��}ȿ�pY�]�d�(�:X�ۖ�V��`���7��+k����O���e�m�T>7@��Եu��̚�x�-�8�}�x�"�݂���sN�\�MҡN-Q+w�����FAN�-��s7�*��u���j�U��!L���#s~Çc=$g��z���߯nN�=�����3�����!Դ�����s��v\{�o���|���;l5���.�:�@�J���C��2�M�bX��g��X8%�G��5$]�i�V���+'�\����y��QO�x�r�V��z�_��d��o��3��#��9`PD�>�;vW+�$�|Mٱ�E�ԥ%��t�(�(π��
�q|���Äұ-��}�5��/ǥ�Ї�71�<�B�:1���e�^��T�Y=J3�՝z�[�QP���?B>#ok-*"�_�t븳|�ͥ���7$�	�$yr����L��G(;���qS3ll��{=N�;P����̢��jt愙u�&�>��f���>9'#o"E0 T�7J��s��2��8
�V3+��K6�� ������|�i�뗡eM����H�0�Y��K�� ��R<R
 ���װL�B��/,%?<{��C��uZ��ݴ���Z�Wc�V�Վqx��h��]�r�D��9H7�����G�fɳ���a
%�ٻl�sD�W#�>�r�K'ʪ7~�E��v�5���2����q�o&��ǖ��|M��e+S����+I�3��CveJ�u�{q�w�^���G�
��|��s�iT|�3"��،�����AR\��������wJF�&�fvo(�b󰑰�1�oC� �l�P�E��o�ۛ6U̦������˥C�.��	��C�E���.1�ךI�z��7�du�x��<bOkF7+L��i?IZ<�w۵��<6��ٚ �R٨�2�ީ��/1���7�[�"�o�� ��֐|'"~�3}i&�^�,�ߜ�۷U,#X.�\�/�8f�����3Si$���px[�C�%2�g�m�Oz3�I���R|�f����@`�޿oƨ�i-c�KŢ�ɞu�	��$�/eu�������ZZ=z,.Xj�ν��F�K݇��w� 	#��9��% )�˭0� �(��,�*�8��/�W�)@�C�X_}����給Ja�'�����5@��)]\��GM��6⪩��*��M[���P�����<��ܐwsh�Ӕ�L s搹�!��y�ch`o�yb;�)J�USp���س�86��y���0e�iW�ζ� ル���PL�}k2SӐ� 7��c�/![\d迱o�I|�D���"�%���<���a�.�̒�-0�g����y�WTę���!�P%�}V�� 2���J��/m�/hN[A�Ù�eٺ�dqQ!���V+��,�1_l�֛�����z�\V�~P<%���>�q� �T��ʝ�D^i	ܝD�G��4S���T~�UEr�տ2-2�PFH��I�R ���[ ��C����� ��K��u^�\�c�hV��	тz{�k�(����_�x���Q��/G���GhL��>:J���C�R [s>�>~4:���D�@EW���|�l� �a~o�]��&:��U���B�u�R%e�	;��1:�C;�Ŷp�v��������N�|�L@A �R�G�����aBeN��/��hj�8�+gBs5��L���`4`�.�(��3:!7���J�t9α���.�Y�'j!�]�	������	vlʰ>�?6d�93��i\���$V��=�̐\�^�v�@U� K"�z��'�
��e@��c$mŖDQ�_�2d��O�[3��	�N���g9�������4���"S_h} Y�h��]j�:U^eU�w�@$q��+)YKz^����r��=�8�~��wJ���#)�M=��Ѭ�<cl�撬عگ[���O��� �0d^~�(?��d;8��QG�� V��Gs�H{���ߏ��d��c�I���Ms��������Ѫ���+r��\;/�~O���DE�^��I=�!"}���Vr?�N��o
�#�$'� Fp�I1qĤ���ѥV��(ל�CB܋�"�%�!�=&+x�i�,A�B�'�t����3����*�����]�!��B�e&����X��yp�>
�նcC����;y8�Dj�o��89Y�z��A��.��
+��9?I�v�����/��%�M��������_�\4��pp L+�/}$Dg]��[�dPRI�A��
I�GI�O[!@����Ņ�.ӳ��w��`4��jI�[��)���C.�_�7l9�G����zc����r��.5d}�8�A���|'2tb�3am��~U�9����ح��c:q�{����;y2H��#T&d�	xzJ\~��[��$�?S�a�ʛo�^hb�9c�W��`��f�����'ߨb$[�*�5�.���Q�~S8F7$��Cu��EpgY�����8�j��ż��G�/M�<f���v��UB���~�f�x*��� ��=Q�\�5�j�u@����?g��4g�ȇAJ��`�{���iȂ�^/�Ȱi����/e@t�Q��Yݲ�N.va��x�暴K��),TVc���R� ^:���%�;=��:��"k��*�9�N��JgZ�)��jW�랆kO;�'�!S��Q.T����+)��	�+bFl�������Rx]K���$F��ԅ����	��� �],#����>|"dO^��LH|�BoYQj3.��Z�cX;���֝Ľ�ɈD&`���h��:���#��9Ơ��b�%��ߑ$�$��0;���>B���V0���B�|J���b��?�����g�KY
1�8��B�O$��K��Q�nI�O���-=�,sG\TNL$I?=��<*��R¶�lN< ��r "�o�+����# ��� )������>��ڳ~�L�$����:?�C*���JOA�-uL5���x�9i<F H��4�m��ͬcO�!t��p5N��ãLq׉O�����[�7&�>���x�E/X�Z%^�]v�Ii|��0;a�,���،RcF	
f*ͦ�+Ŷ>)�y&,p��&52h�����SG1L��O���c-�����b��r��,W���j��@"y�b.P.�������7C͉�jW_j(�v��E�T�p���;ߞ·i1瓞��Jn�ܯ�a9Y/w��j\��[���7���_W�Q�3���S���w(�����S�:�¸�|]�A6���k�*�wņ��,�x�.�,i�u�14JV��D=湚@ӱ��nc�)ve�ڢ��l�����dWV�m�0,/���e��A�w�w��C-_�aA`��J��Vе�a �/�����T(�~�w{�: ��yOm���oS(��]u�7Ay�b��������L�s���r�*l�׃�Jpm?�9	�A�/��BQq��O���%[z�宓{�̛�hF��H!�6普Z�ޚ�+����-<C��+��I�zV�X?�1��ǝ.��!���;�>e���f��ӆ���O� ����G~Cǵ��.�{�@G�w��Z�t�&g�&o�9_E�z��!��A�{��<�� d������^��T��IZR��
'�T��/�-u�_��$��	�,�L��2��|�0{'��!z�:�piܔ�C�s�y�q��%���_@�����g��dȳnZ�>A��Z�(Al`[o���b�>{|'0B'9�X}�rV@��!b��uDLG�[�U%^Yi���Ib��J 9���-r����?���8�}-�� ,�R��;���`S:�I�$���04���7�?ￖ����'ɝ���r����Z��
��u����{�%F<m�|f�X^B�N��\��D o�t�[�$��l��<�!������k	�Y�'j)���9tqa�Z��A��bЩ�u����c)�$�U`�8�tخ9)����0�{2D��5�) �����ݛ�rk�*5���&ȴ`�x����X�e9[�m�h�;��}ǲ��/���\
�fb\]} w��cA�&�W��D&s�'�<P�`ȅ���d��	�.�*s'�j���O"�C�jb)�����`-�]�}�N@�<�X�*�����:k�6Ѱ;�d�kF�V��_��mD���~+�6�תd�;�6=���ۡU�38|�Ķ����ksh���j*�|4��t�Bu�?ch��C�ݾ�'{D����=_4<;,3����mj�N��ƃ��� #�J��v`уԖ:1x��d����*���R�]����{Os�P'b�R�G��o�A>�%�Ϩr �{2�V?
ʏ�]�|M�7:�"I��	S��E�&hH�b�Y2�:O+C���Iu�OCo%�����[z�i�1g��,�M:j�[�f�[X./��MY!Mw�R,���%x�}Zx��M~1S����=F�z]#���a��j�����C�t޻;��#����<%���I0��v�]��	C�����jn��<��mX �2I�.z9WQ3Ut���d�@ϱV�m�~V�ń���WV�p�s,2|��|x3	�m�-E��r�u��!,�$11H41�� �[�*���}c��C��L+���iYp�2��'J}@p��KMv�3Ys��$}�*|9�[;!�o��)�����?Z�˾�N썑C��<0��,b|K'ۙEȲ]�p�m�]�*·��p�����XQ ��%�y��:���`
�^j��=
$5x�QY�����3[��ff�Ȧ9Er����IGೇ��W䥍!�Wt%߅��.*��j3p%\�ukϨ����R.: �p:�����蝆[���M-�"������Q���p}wF�a���% �L�݀
w���s�O9��x2�K�9��N�]>Ep�mH��i[�U�ר���tX7��m��< ��O���~L,Z�S�q}��4�?'�bـ����հ�9p��� ����0�{�f���������Ū�_[L�	R�D���f޻�>P��){x8���<%�'űu豒q�������m�z[Qi�������S���}>�W �:P6��#�X�G�Kib���C�� �;�JO��>k����{C�wC
�U�H���@2!
C�Ib~2���Ev�̤�:����b�A��\v����K�Wx�اU ��d��d�>Y���o��42����-�U ���~�t�N:]A���qvuO��n2G�ة\q������
��Ɂc������'�����D�/o�Gk8��}7q;�xAi*��V�ld]$�ȁ�8,p|w~���!X�%���*��_��V�+��Z&�'L��[xs[>ΞM������9��<��	��`�� n+����6ʵc��i��v��}"]��~@A�� `8�y&�禞�~Q��^��-<b"���&���U���r(w���c{t4�H���n|V�@�̐���4 .��LLJ����c����9d~M�C9B!�3��cEI�[92I��6*6+�Q�Q�����h��n��J��-���`E�q�ܝ���r��XJK�]�K�.��rQ%��u�kS�p����XSÔ��m�u�7�l�?��`x�g�?b$�>��.gʍ_���{��,����e��vn��>�o +��
yf�霢8�����f3��o �yK���P��X�M�{�nt�|�f����Q�ryNNŮ���Ǜ�{&�0���*��,��t�`�-��� �@E��L�����p�T"�&��=󪘰������w��F�鳤�c�#����na���$�n��x?���l��F����q����u��%�F�c���䀒W<�} �\?���Uȶ��r.�2���E98���0>҄.�:k� "�����1��j��1�����΍!�"N��+%m�dO����bh������H��,�M�B�cRj���}��򉴼�p�	���\��;�=tY#�צ�6CZ��V�_��{7����*�)f7<3�:�5;ơ��9 �Q��l	<�.hw�Ŧ����hp�o�.�[����Ÿ��\�~���1�">����n2|�F\{^��h���N�p�0�x���ҫ�10&SX_(����!�lS��&A�p/LCq�g�%�,#o�c�l��$�sxH]5/���o��t���=�l�w��3N��D�{�5T�5�@mLV(�Xh=-�Z�N�2�z��Wҹ����#$��7��Ea��#��}B�l��\P��Cta>�ǘ�^�\Z�&^k��=�\�߈(6yr2qz݅����(�B��K>4pa��N��=���--�ˡ��˻�L3L8�%�G��l�gY�!ц�R���e�
+�q8�BV�@��_�k�o�X��~�^��>rֱ}j<<_�T�9�9���N�:e�����o�L ���~�i]�UR�bQ�8J���ђ�n3����+�8)�{�%]�sq��w_=m+bMc瑴�6��W����Y�X�<b��D�J@j�WP'�+0M������@�GqN�U�[���f)5�����l�c��=���@L#���Axs�/soRA��+ˎ~�{ ���&���<:�|���\r�p��T6شc�׽��p��i�&�j�4G/Q�.��Z�+�����#�����m�ݪ�R�|0��k�AZYZ�Ȩ�<��S��hO�%Fȩ��TN���Z-�k���(-ш����a%U����X�-��l�̐sI�pi�L	b�\��R�ۏ�r6��k5=]�F��pp{�d�k�噬b��鵄w�W_�~�=A�ɮQ5d��z�t�9'��^Ϭ��7 WuC�⽟ ��>9���Nb`�He��J0�@Bc��%����xmkm[�W+��N�V�n���6�p��2e<8�Dqǃ�DSo������P�.+�4Ӂ�`+@$���]\�?;�J�h�?Ww�PG�?�}�km%���~�G��^��]ڄ�!Li�����������H��|`�h�tq�
���u7�r�[ֵ�T���13�ʹ� ��*��AV�2k��_��(h9�
IJ����N,Y�{h��g�l��e�y�'Q`���u(V����|n�+e��|�0>{�ԣI0I���A"�_Њ�۸ ��� ���'NN��2jO`URM!'辗���r�Sj�Kp�7:AYcA_�7di3�j;��J�h�0�@ly�n֣�/�.Y46c�%�	-$����M����	�4�׃IΤz����##ea	�3klѻ��9���~7�> ��f�rع�z�%#r�ࠜ���:�C�ɶ��M�<�� �Z)&�*��5t3�����?L !�~)��Y�? ���p�&���ݱ�4-6�1��d��FW��'��Y�u�r�fq7�O�f�T��֠���q鵞g�x]��Y���W��b�yL��L��=0���o��W ��?�~���ex�8ȯ��� y`z&A��Ϡ����1Ό�w�����y����'M�J��xr��*��c��X��d܈���;�K|�T���g�o��	���##8����Kc8��E���0�xB�����k���k�%��y0#�#]睙�����Vr6�h�:�5��꘽ͻ�9�i���`�~2��
��$W��AO<�"��O@cʴ.z�x��G�p_.H���Դ�����`!�ڊ=U�.�t�W�G׽���C����Ҩ���,�m��-v	�MM)霴�Q	��;}\0V4��c�M�� V4��iGL�n�BT���{%�SY���muQ��{�@��*t�_��nO�V���2�Ue��Y�5�R�k)�C*�=�Ph�	�fD�6({aË���h�X\O�ţ�T�-�T/�Qņ� �V��0�t<�LA�TQVD:����2����ɀ��$6Z#}�hLzt���X�@�}7���*�ν�J����(b��L0ǧ���|���i	qR��J��C�;U}�#�Cx�B �t��f�#O9?�탥?5N/�uO\�UuZZ9����wJ��Í#��?䬗��}e�U�Pz�"8缡lF�.��Ƅ�>��b�Q%V�״hc���adU���Nw"̟�AT9M$������@��ҿ�~���K�p�#&�]Ƹ,PaH��%+��
��J֮��� �׆u�Ȗ�)��*��*C�`�e���vW��>#�=�S�t�l�*������>^9ۄ��Ã��	��O�J�b�����a�I6�&;�Tw�t}ik��V�p�mH�h=1k�6{���&Ha����U�����|H����uƮ:G�6��Og���!�S�o�1���<�+��,�@,�Г����Zaόo�m�_�.evL��{��T=�]���ʇ��aSP]e����gƜZ.Um.�坲�!�c��D���jO��*aC�]cÉ�/A�v�*��UkY^���<�5��%h�qh�fl��k�n����+����y���	���ہ��0�2[��l��}�4��g:��- �$�2,ѭ��sd=~��8��[3k�q��	�fS�h�Aqp����2�7�s~BCa�N\v���`+ǡ��ê��;I�^����v�)6���5k07y����8N��Q|��Q� ��.��0܋E�Q��Y�CX�:K_���9<>�)��Uf�M���BvQ�F�t�7��	�K��:���)�}���f�,�LT���B?0���{x���	�z/��q�&X ���A���tW>zk�΢�W{*p�_8�J�w�"qђ�R� eZom���1.�Y�/�6[qol�	�o�Ė��v��e�V6`���bd�mS�&��f�������٣�f��9�7OL��`۝����[��A�
��o�P��U'��.8-[��W�4/���
R"�3�Z��ȗR������+�.N)��-r�/ƹ(fZ;��s	�i.�%�c:2YM��>F%��1.�C�/PP1M`�_��&�#)Rl4�GP4��RK<�M��.Kv��{�_����^�
���wW��q���������q�kJ�[���<D���;�}�eG�Z2��EkJzv=t��}�K+���ZG�z���Ƒ�.�]�#���9-Y�v	��}����A3���nZ���-���ܓF�����*���'%�yu1�3k����|t���Ksmv�hKJ��I�|h�RU厡0]�vm�L�hn"��ɏ���-Wn��]a�:�L�VJ(G��S�;��I�#)6����/ֲ�/��b,��	��T�� ��}�Տ�.�1�2|�i�`�"�b[αM�*��PԂ0-��)��KTz��7�,��ё�6��|{���1Yԋ ���F��!�>P��~�Qb�_��1Jx!{���c���H[��ȓ��g�q6�(����q��m^�-DU;���!�U��x�{j�����Ul��Y�T�8e��	�E�� ���N���٧*�ƾ����*�oC�w�g"B��~��ò5ۿG�7�C�=��Ucu6�-��+��)'������&� Y���wkf7p�mc���zĴ5�=)�H\�Ќ�X �,BuS����u���7�Y�X�R��0M�VFa�O�T��h���TèK���7�au�;,��X�@��^��o␍��7C�}��'����PF/���k�����3X����L)9�n6��S�<�]����V��X���V[q�,��L�悝A�[1� �)ҠG#��C�-��b�:����?CY�GN�u�����
t�n���Ʒ*`�i8p��x�o��c#;#�B�!�����Г3"�H_�ѹ�"
� � ���(��L��V`$��J(����)��[I��y�(Q�'�KL��Q���ʷS�����"�Y}z��"iD%gY<��z{���=�&�6�laH�_K�1洑ޑ�R}\�S��F��|�����Y&MslJɇ x7�!�>J.��@;g��lLx�뗮#��S�p�C}�ɐ�M_9���l����z������>�����O?��{B��߮�mv�͉�M`/-Ȑ�C�{lk���h�}���Q�*T~O��1I�ˮ��q�hIZ���x\�khMa�{҇ɫ��9�*w_<f�mt+�V(�����i�\��m�A?��O0eא��˂�_��V�C��9&�h&o�P�M���;JAV4/uI@?��$�4l���PN��O�����lL��õ�o���H���^Q'��
�b�^��j��\iԮ%c����9I�b;A��p\�'WA(�$�����T�<!���#���v�6�	�5=Z�h$���7�f��������#�g�O���ҷ��P ��A(͞�|MCnf[�n2�p��a��l�Zm���oX�ZUM�r���\�Ԟ�l��EN�����_3��Qt��dP[E:5`��m���m���Dx�?P��v@ �ed�7�J3P^|lrH6+j�G�$�mpR��,��Z�&K%ω̃��w��`��M/7�a��z��IIBr�2��4_�5k?:�1��b�J�̣��!iG��l!�m���|%$e*H"E݉������Е�F�:���oBT%	�K�
J�M�'d� ��	@��O@�+��>ƃ��h]FR�Ҳq��rRA��&���F ���=�CcW>0�X�x�@	�P��|?�g�m-v;���'���h��q=P`lK��tgy?�niOo[�%�o�S�X����g���J���%�`�8h�hv1��	���1׸�EWN_��˦F襦Ϊ��m�L.�$��z���L� 1h����`�mnB� ��SUʌC	�t��`�A��Q|ʧ�R,��8e?~��a[���U�O��]�9�HB��G̊�k�|��_��LG��ͮ��r<��
��Z	zD�r:<�}�R@�#b����u�E��z��4ua%cr�S��'��W!B�Ez�H��,w�����;�����i���
���۰p��3H�����+�~ҁ��\A�p��F���?��0�ջ�[�Q�Я����yVG�O�95\=G�~�6@�,�4A��TænU���kG�ON�����lYrC�^���z;���yi	9+`9����n�`�~C�%RTm�-5(a���Fx�k<?2��t4���`�jQP\l�8��N�#�GǄ��b/�x�;ϔ־��X��kN� ��23T޶���Q�
���Ď�	B�*!F����R2�>g�k��_�k�HS�2��';�T:�i�����(\�&c��!�A�!��uʀm�$����ЂA�Ś�bA����������Cu/ܫ��~��桲��Յ��@�!|��{_���� �X'x�$u�P?W���HI��D��eWR�|�Ғ(���O
����y�/��N̸�1o��6e'�������+Ov���R��p�0*)Ǳ,���j+����ˎ��{�:*Ns$������Ȱ��pY�)�a&A���n���|���:Z��0B�0Q����x8t�Q�)�M�������1�>5�4f�� ܑW����u�;���ā�@�� ��d�դlĆX��*U����7^����}0���4��TE�E�q��I���B�9�	óBܜ����wk������ȍa`#tv�&�^�C0�@Iz8i�Ǌ#�&���b�3�y����8B1�\؏����X+Ɯ�D��Vb=.Xp��6�|�I����6��8� ��z5���f�v� �`1Z�PXxb�g�He�mp�$�R��_�6�C�wh�ظ~�i���^�H�]Ua����{��6�?D�L�[y`0�,"�X_��I��ql�n�>�sb��0}�a<ݞYś�!��/H�m�nº��?^��������S�{׭޶?0z���I+X����������Z]#�|��IU���p���*�&+�������7��M ِO^� ~7��p�d����l���~�w��^c��&�YD:$NG��Ʊ�V=D���"��-U��>��]o�厬���=��r��ú�[m\�j���'�s��{U������uUi�ʎD`��Ys|��-�6���|C=�՟l������E�l@��ʿ��?ۥ"V������y8���x+-I�N�O�D��BJ.q3F��=�X�IPE��|��O� ֤��"��6S�?�!�v���Q�آ�Q횭E���b<u�(�v���u�F�/�0I��Vyi���B�����3�������������~�_�	ZH�K���a
�p��,jF/D�[_�Ea��ն�%0:���k:sC`���!���9�<��t���	����E�܈�[��: �Nf�����sO�	-(����ͱ����p������ZO?�Ч|���Dl���[K�������B3=6�K�R�,}\�=�:I�x!m�� Rp>�������ܠ���'�H���Ӌ�[z T�dv#	V,	,�tD:���z-�(���z�_��$�A�8��>��woZ�;�lƑq��fCV2o0�Ҿ<܆�p��&���X�8W8�	S��đ$*rϾ�a~_��6��:�j;BO� �,�E��q��ߡ!\S��u~26|�E���k��F��/M�s��R^����k����_����`�h���4���[���w߸�[Sԣ�*�����l�/E�;C�
���������	��A�==���U}Aː�i�	��qEJ���b}�}��_�c���d�W}�l���R9��r](��"��?��sֲ,�b��nʗ������]�c�6Q�T��5P6�[А��%C�h�gŒ<�8ՙ�H�'�h�������2��@�bR>�@�X����i��~B�R�˞��{G�UA���ĺr^�*<�|T������w�A5-1�Nc/7<�Q��-����U�w��܀+��<ϙ�N=i�X�yZZ�͟�c�D��@�fa��\�����ї<MHz7Q�v�ӳ�8�M
�F��e2Sȏ�P�|��)*Ν�h(���Z�f�@jn�΃Fc_FX�� .�Ԝ)�����,4)�1b8q�ʿ��qٲ�ZMd����,��=�ۼ��E?�V������R��g~����wB��5�&�#?Һ�5��#�cb����Ґk*�o�0y�-��S�Zҭ�-��H��~ m�·5)�=�P�~�@@�Q��<w,5��t��L�|�W�8�}K�5��q�&�(?�p���0\��l�q�$"d-�Mg�i�����[�=)��pN��f��	e3���z����3��@!��T�8�Q�]�*���4�ߓ��?('M �ww�	�R�mV�4�;q�1����Xj&���=x���Ӽ]T�\
�gqw�X���5�$���V��B��o�ʌX<YCsm��ĭO���e��iź]�f�]pJ�f��=��ěw߻�҃���r؄��0�%��v�� UJ����e?X�h�1��κ 1�/��;�'��O��@ڴJ�?m��^j�f��)oO)���wykݣ�Fl:��/HW�����n����C��*��7m]&E:z�qh#����=,]�n<T^�|_�d�X���t�� �lO�$�W�(����+��7d�%�6��88�}v?6�����+z�� t����$��h#���t�T�8�b�.�����g3'fl��.��Df���%�G:�z�ד�"�q�1�SvJ��w��[l��GݮV���ޚ�쫤O��M��V渫um}4h�a`�0��~�1�dM�F�s��Р:\���8��U���w	i�(�����[����%a����v4�]2��µ�l���}��)��Dp��e<䇼o����ը<�}u����Du��;��=�^MKl�F�P�۔����Ͽ�TN�D�Z�N�3�/�K'��>M�U��o���'h���������&�֗��W�稨1��5�=�(�D�E�r��)~���Y^y�y�����Ĕ�Z�/1�t)��T������62L��]�Y-E�)�U�Cn�r��t:�|�&R �������t����$z�b�r��&�٘�!��Ǭ���<M]LTy˝�l�64v����Ի��4ǭf��!�/Y�n�8Q������6��4��n�[*5�	�+.��g-�<�j}�'�����D^^�ߪ���TX�������WFKciP'�^����K �H_�QM��b������*�JRh���~�*�hO�����C=y�L��_��{>"��m��\�ǅf�?�h0��X�]���( Ŷq�}�I�����I٣FK%-˨m8�!���ێyo��WS3	��J�	�����\�������wEF�R��@��.A��t��Tjp'�k�:b�/v�z�K��9��6����\uh����Ӫ��➹7�:q>5�\õ��f� �$���ݯi��jD�tFMm)�V��!�2���{(Ig�Su���	�xE�$\ǧWzv�|ԉ���#���om����� ��z�hq[�����+y{s E�n״�V����91�՟;p=��
��ҏ��}�����anw[��F<��C��kJ��	�����<p�OE�V�A=���yh����ν�~�Ȼ�Hܸ�#d�ߣb�#+%����vՑ��>�H���v���A�-���+BM�X�/f���}��_]��@�T����)��0	�����K�\��*QV�<y��3^L;{���۳��t�\ŏd�}*	�6�QӼqA�W���X9zJe��z.�滾]ɑ�b��J�M���r1'�*Ja!��Rd�-�(ɫ��D���s��\_�e7�s�ߓ!��A
y�Os��
��b"�ab�`�d�P�a���@M�Î?�R�!�,�R�Ύ��$�!�K���Sc�F?أ�ѦF$U��{Y� ܣ6K�f��h!B]�kp`g3�@'G��Ȋ/Xt��s]��X]��KYB|c��Q:m����Q�\�뉍�>ZB����o��r7���l�`͢	�����Q7y����bq`�$�E
	���6%����������iȘ&
``c�!O��M}4�6#U6�
��L@yu2��:�]�G����S��c��u&����A��׍��zU5e��C���m��i�D�+����f�]�L�h�K�9"G��� ?n뱜G�1�B�o�0�NSKxC�2G��j9���`������}�;�2x���� ���|���g:�'xy�OK5O�����_ &�&o�N�K�#��(r�������+b6�JK����/��+�< 77�S�d)�l5��mB�����؋@5�(����q'%a��ټ���lw���V[0s�pC��~�TUA�F��F���ݍ7jW.	句+}����z�_�x�Y��X��5��Cr~��r���J/����0cM�t����Xc�0���PPZՙ�e�(F<��Kl���6,WA�`�����r<�YA�/c��c�l)�L��H��o+,<��)���V�?���$E���v����+H�B9l��Z$�R�σ��e7(g��������=�����E]`�W��`O��ߒ�~ʖ�����C�l�g�b�;�����˹b��ї���З���2x�يiZ���F�(�r��k��R'�rv9�3��Z�j��u�+(��X�/8�G��FPb���Å��5���c��XA�L�
93Y�Q����QWV�y����s*��X�ve��6�!-��[RX��2֨�1�/1�H�Ն��޿��!	-X�n�������W�)�\���c*��W�3�=&��1��C�l��z�������w��j�j��$�-�~7e)�9�Ro����5�D*,�&�g���}��"=y�K�;�u����>n�|Z�_/(���a�k�sw���S�vg��	0(�0�	ȣU:�uJ0!:Cm�j�6�΢�OMAt_�wg/yX��\�bet�B�{�]`�8Q@'�c3U�^պ�(�O+���������^�r:���L���͉;&�.$�!d���!kK�R"�򱑫��t��(5��^���n���u^��Z��Aۢ�xE��2`�0�"Q89��5C�4�f��ŕ�y�;X+CXw��a����)0�[F�W+2Kb:��̍�0͑ ǧ��{���Z�&��g61X��/��� �FP[��Y�3���a��}�\`�,Qo�)�����:��^n��.nZ-	���zy��AG��PH�-�D��Xo�ݿ?�@e�)�/�o�qۧ�O^�Z%B�:�2
I�.s��b�DY�U��������'z�b��U�(����&D-�L�P#�jC.ie��L�_:庫&4D]�U7��K�H��Z�����ȗ���Fs@�a)��a��ZU��;#*i�RV�E
P[�~*��'� d/,;���()i�`�E�V�H�Vb���L�`۾��_��z\%�1��U�� �(<���<Q k���ְs&���i����Z��n���IO����B~hm�-�-v�����LV�ս��D0>����z���^EÇ۱���e��������d6߽��p��zpu�I
n�����h��ic��ÆC�m2��c� ��"K�!���ҁ�w�4}�I���	�r$� ��NW��! �DJM���7���I�6��/�ƌ�gO�i�F��D�d�\��c��^��픳/��I/�����N�(_����.9Sd"T�}B����x��ʢ����f�L,r+� ��(�پ�RZX)�+�X��݂��ܿib���w���Pl���6JI/�n�A��v�3��*Y|�eL���Ⴛ�VV�6���jݐ��	�����(���z���+u�PERʔ�%N�A���:5�땫;��U^R6�ok�3��ĉM^�$eqq&�	\��Ek�C�Įc���,P�K���Rď��-4��n����f� ?)�����hǑ�Ü���uǼɀ⦌/��،�NOi?�xᐅ9����<>i�[W���'���|��v���aп���ǋ��6�S����u��:|b�^#�197&�9��v�K�4�}i�#��H�pgq�˵l�����及�ڋq���a���O��
U35�1�d�Ca��q���e�7�:�k��;�i�_�Z�6��������a��E�8�n�A�L$�a��-���6o�PņF��M�JY"d��$�`U,Pli)�o��N�Q"�"t�����uk�
N��Y�(�
@{|:g����ʆ�1h�8����^<�����N�v,�Ic���g����Q+�j~RʣEg�¤��R��u���J�^IV�P�[�qAt_[q|�3|馥��G��� -��Ҟg_ϭߜ���%�X�۳n�x�NF�=�(���1V���z�ٓS�t8��̎�)Ɉۼib1������*U�yes���i�=\�Ko+~�ܼ��k��n����V#)��	ES-U���/-���L��
*9� ���C��Ű8�iY��L�X6��ʝ�ݫ^!��f��H�KHIuq<)'���R����g����a��ѧ��\����G\q�52��NRu���tȱ�u_3L����	����Ԏ�=���x�ʪ|���-XZ��</��2Ã�c4�[����\��m�)�bm~]�~)��೷P�IK�T�̩�l��,x���f�{��1�KH�^�?��8�5�ϱ?M'ckY{�6�s�ld��'�D�4��0��BE���*N���ߢ�ܺE�Zc�
����t�0e1*q������,��9֔聳ʐ'�NH��A4�W;���O�l����Df��|l�g��i\@پ���<2E���+�s9�_��&.ِ%u0����*�\|�#��ׇ{���ف��֗�6�|�:��r���(h��Dӊ33���Y�����ޱ媮�M�̬XvL�wS�8�4�W��͂ҸY��
GZ�B��9{qy������(���pH݋��0}��.�߲�rw��Z�ĝ�o#,�X�"��-,wʽ?_+{�X�tV�
���F*�+ߋ龋�'�=ygD^#Q� ��j��w�����tH6���5۰A��®��7f� =t1��r5���B�F��"(3����tN4� ��=������o�DB�y!]V��YH���(���T6,�θ��gv	*,pTS�5L�G�	��X�}�Q��_�B��>P��)@��ୀ�P���։^��I:�F�E�;Γ�x{�Xl-�"dt�u"Pm��9�G���m��7��_y���=��%,uw��[�!�8�۽�_���b��qz���4�eX`2��khD��ʴ����ɳޟ|՜5:��c�`Uu�;�e
_��n�%��9�A��F͙�2\�p�������uI�c��t?S;}�(`���:�%D���ZcS�{�yW�R�Q�����uG=�=��W@���`�/��_��lCIH�#��|�dcyM�:1I�>n����C�R�����-�z1��P[$�d�uBSI�����=��#iQV���Z�¦xO* ��e��u��Σ{�m]E��f��#��D`7�I-?1O�2f�li�/���Kf�����Q�6�O�%�8p^\fl�]��é���n4��}`6ZbU��~`��y( �|�l�d]��im��hV�L��_�U��S9���,�"5"�6��Z-�8$,�vi�Ӵ.eU��W0Gl?�9��~�6v.j��� h�z֠��S�z�Ų���%�	@J�+�/e��<k\;@i<���)��}�X-ŗ�G�:��P�����C�JX#����(�i��#��#��F�Gi@�}�Q���}�+��1��i׺h�3�9��^Vf��a71ƪ�-`�����~?�XU�9F%&S*�R/�;W^��%���%��n��z�GD��]�^h�����'��0��0Ew܉ ]���}3�!����i���2!�o�j�H�0��(D\h�Y�|0b,'ƺQF<F���Kb���L?�;��0��nC0���kMՍ��$��Dz�o�)^�1XA"���E:@����� ���*dg��jhjB�
������L��UA���/������MG����M]����+�>�u�����Z��]t>��̡�Irֶ�w�d�E��D��l,HS��)ʭ+��^��6���R1�!(d�H����Â��d"��֍Jke`a?>=�8	���6�NR�1éyC�?*��Y�:�O7�me�S�i�<�e�`%��܂�Ù����[��3���^��ԩ�GD�CN�:B�=(e=���[������k��|��.�!��R���]l'����dHɷ��\�{���|bK�����y! �@3�l"��H�tN蕴����v
]�V���|ۉ��#E?��������1�0`�*(��B�f�y5�v�4��?6'��Èq�A��~G�@T��a��L"�躘<�ĺ�Y�\ԕ�΂Ic��nr@l�u7��.>��5���k9�i�������M8� #$}/��k�;o����g�����'��!�)�?��'�:�G����Z�����m_"�ꘖ�5�X���Z�]��I�mP�Tܺ���t�hj������dh��!&�՝c�����B%y��8B��{�p�Ģ�Q�_֥?<���".g�逹��\AH*T�L�d)�P-����/��Zٱ`�����_���Y�xw�$2��BUu���K	p�l�j2Y!$�.�x�e9�~��F,-��|��W�A�Q�I|U��/�t4w������F��a����fomJU���gd6㢟N�mK{��:k�T�n')kuu-O3�f��M�ń��'&G��R��2T
r�G����4�;ؒ�^K�8�9����D�X������[Č8˙�����qM)�v���`h�t�C���i�����s68<� �-"�*>s�\Bm�Z��0&�
&��-��e�O(O��а�a�+�1��G�ה���4`n�]i��u���9�#�k�/�l�����2V�g��d��T�o���&(�Y@=X:��;wW�����Q|��2��nX��|Ŏ=s�\@�&N��t�¼�ŗ���W�����[��՜šM��Y�ɩ� J�w]��;�3�����@�����9��;a�%'�l�P���D��ס�8��aG�H�Q~n���x����V����v1/R&�W����?B�'����m�:^�+[y��������G�->}D8��֌��EU���q;���v���j&i,��.�#}Y�M	�l0D��ϼ�X�d�Y^Ɣ%��K'2dԃ%�L��䮏��i翈Y�=����}|=��L1{�Ȓ���H�_4�U����m}�/i��@���sUt�����dO7��bX�{dM����`��:1&��{, ���Ӕxz~��"<�V�O�`1���,.2Y���	�)u�0�'l���}���gO;߃>�E;�� Y�~��F��l�=��BP�u�{9�q7c�9!��"̌bΞHB[s9�7�������I���K���ϵ3�th`p@�u�*���:ã��A��N0 d`{O���`��T��T��,��q�2�:�|B��v������Nm������D��k쨾.K��\���r1����Pڹ�$ա�?��g�77�E��;���HՍ1�%��C;��#U�508�&�쑹;��nWP�v1��ǚ����g���v#��$ͳ��Z�T��O�V�1K��7���n\W��!���J k�gx�C�����51�Zx�Ӗ�b�]���r��`K�UK7�#U����jv���#�ij(a5�7!I��+-x�-��f:t������Vl�*�$�YꀫLN������p�H���E�9���\|7!{�fx��B�w�|�Y~I��Pߡ��U�e�m���EV����������5�e$��cz�˱����fY�ƬYh��R�b;��1�($�<������1l�o�e�A�\��y���ǈۈ��s������T��4ڽW�٣��� �0ԄVƸ}�M+��o���@� �F��x�ގ��CLpa����Q�w�~��� ]$Z���$�n�u23�
��
��iɎ�{{���[�,����#D�X��<��p]���s�WZ�d]u��u%b�bU�&�q����6�2�>����Zo&.
� ���^���Ef��ә8�s�3-1�"e��
Sh|V4����,}�d����*��Ay�B�/�m_=E�8��7��nep�ی"�*~�J!Y=�D
=�@#�K�xo��`pd�h�������DJ��͕g�`��
�r�E��p�u��N�U ҈{�+�DӉg|�`�BL�(om|�P���_����#1����͝]C[&��{��k��cQ񝾒ڴǧ$���%����&�l��H�_o�LLf�����v{���RC4�H���D��V���|�&EUU��lh��������Aŉ�^�[G'�@#����5�n6-y$/b{G��T�.�j0��{F��X����d�x>���z��Ns����cﻷ�Y�_#TUg��f��ZPu�pG�J�82�T�]�����ƻ"'m��T@Н8+��Lz�V���쮵hzw�C%���s����9���mT�{nQ�v�,e�uX�QT�	}��8��(�TԾ��Ԁʅ_\>��'↑�t_������½b�YBf��m����l'�v9V
�0vg3#�7����q����LŠ9�z�D`��B@��6����w�[.LՎ�@�\�#nr�'R��@}U��>5�j�0�a�	j�XI$����@3	ܑ��H�<�@�і�Gx�W�m���%Sk~�c�s ^��,���n�@�zQX(h�u��Xs^�y6����p�)�{Iid��Q����	�pB�`=2Up�]���1������z-�Y�W/#*��b�Y���j�˓`ޮ1�L׵/?ph�w�ytj%"Q��f�I�6�E<��ŕE��*#�y�^���>�.4q��־�x|_Kwld��1�e�Op"�$:����[�G��E����o�%'��f� kϼ�*�DOr��*�o'��מ9���]�>LoQ;9�(��������WN���Ť��m�N���,6wp���k]��!�*oP���gB� =2��f��J��e�{�[M,���pr�Ԯ��������V:��ߟ&�yv�J��l�NͰ��p;#G�����I���}��Q�/zN����G{E&��Tu�
!C���%`�B���9�T��̜λ�)$ٿ~���9�q���w��I��^��<�ޟ�H
-�1g���Ҋ��j�+�o�^��y�z_'
F�E\����%�;�Rb-f�߶�l7��(�� �	�W"-�6:*躉�g�5D�o���R`��"�&\��J���8�:3�w_��Nт'�qh��G�-:iY�nF�M�+Z�F�z;�c�2[U�/I�D���c�f9��XI�>�|l��m;�_��%GBʁb>�����V���R��u[P�n��<,^s��&[�<����5�z�y��I���^ g�(�#6}s������xq��H]q�H��fYs_p~���9͠ݬ��@��Q�6/\)�LC%��j�*򳽠��i���˟����`Ϡ�c��*��5iF|gf��&).K~y��Y����9DW��W��]R�zp�l튰����[7����5cث����R�������9���|v��oZ��<��v������Ԏ�1R�1���>TҎO�*�:�Y�'#_E0(��zX��*\V&U��ެh�?&������	�n)vc��f&��}�>�D�auv�^I}K;�W�o�r�0m�f���췮]B�;	��,8�ڟ'��U�S�7U��1�:N���|�����x�,&ل���N�K�3p|�<4�^�3�������eਕ��媷��K�7�.� z�y�)�����_��9�]�݁Viop�[��n�C��mVi���v���M��� $P���۞�q������9�@�z	���|<ཅ�'\Y�-i@ϸ��{�Th�}*J&�L2�G����N��H�|�?i�U�������țA2>O�\:\:�%�/�b��d�\nCE�h.dy��$�!����s��^6^T�4�.|�?��J�Y4E3$̛�)B�ێ޾�W�Q��d��͘�+��˭rz��3M�ƶT����9���-J��|YM��*2��3�kE���	�n����f��R�.#��-a�ܪ����/N��ܹ���� �j�I��[�{��9 �c�+$ܲ	Rz�MN�Q2T���O3���~��/�����屬90 
&�R&6�W�A�� ��/
��C#�����H�x�O�� N^�W���K��},b�pm�W�c��PM8#�2���WP�J�)��[{��w�{�5�� "L>����!��vhM��'�
B�D|P��4�{���ˆ��ަ�3g�:�-�_A�Z��qW�DY��vu^P3r���d�џ}�A���Z��^ɝĕ ��8�s:���?��%3���0�	�):V��:5ֻw5�}����;/�����!� 76S�{01���,6�ۼ�vǍ(Cޝ2$0X:�4uЩA���,b�8��b9~��wX*�?��a��rʠXׄ`pdl�Ӳ;������i�el!/�_�X<�@�h\G�)�z�!g�-���:�ȫU�g_{x���i�p�H�?����(G�m�]�F�%�ny�� ��������p��N�m�C��hT0�c�&�G;~�6��~w޶��y�Es�����H�^;�ӴI�iT N����M��'�TK������UY4�ը#Gw51U���ϐ!���W���C,,�,�tUϳ$r�6Ӻ�cq�+V����l򝴇~��u��{_*�dKg<LJ�c\+� .��H;�]/����v=8�}k�����U}����}��$Ђ�:D�� �׹�{��
����L5�i���c���ղ?k�K�̹H1p�)b'.R��=Ƞ^�mDv�*�O2Rp�r�գ��i�F�_�|�������w�2���H�^ >ѣ6�Tɱ	l�XM��=�x~ F۴�~Y��ګ^a7��r�� >Dk�$QI� �c#�c�}2���2Շp_�#�Zu���/#[�٤�����3����/�/�r��.��&gI(GVqb�tB�EǤ�6>�cv�K����?���g��|	�1������IÃ���P���n	]͋��gU�8��o��.S`su�@R���+��wE��râw���q;/o�a؏h�5aI�a5���N=���W�\�ɝ��ު�uX�(�?z��4����O~F���� ��5�Dk@��`�[|gc�Nϩ��G��.�5��h�w(�TB)!�Y��$ʞd�tT��h�R�����EW����t�A��xtM�a�k��z��Xq9,�vD��e��3W~5��G<���(D:&h�O�}o�?$��6
5>�Cct��R�(}�I�D�������ē�P��rpZ���^��!�R���׆rS4�
8�w�E|TP�C�7N�������~ȡ�'#�C�<���4��d�R��JWKC�4�h��~\�j������/sO�Q�o!A�-���?��{+`���.�|��,C�IP7��kv��)��#��a��!��Nh�����y,#�$RBU��%B�e<���A�@O9�8�dn���Ѐ��XA���3p^�&�$cw�M�Z'����8�V�5�����v��:�ͷ�'�')����Pɒ@\���Y���.׏�0��n��A�"��

��?�q��CN��q�z=��n�P��)���.^?V�F��ɲؙ�����I��h�%B���7]8�l�������CӀ#���$�^���q���t�#�d9��zq�k3 x��D� � �S]0m�@�9%��8Ё�X�K"��2J���\"$�L
y�T��
|V�!U�s,bzJ'�z�1R�zw��a,&�����SuѯWtа��R�s#86�j4<�������ecO�l;q.ǎ���#�a.d�V0�Q��3 Qk���:ڜ�1�bH��p����M��U����l�	��!� �mJ.#ۏ��㽾Ͷ��C88�bۉ���&I��bt&�_�u�8���ͯ�g_�%�)��T{I'<ڕ"�G�=�>e��c��-��m�����M�9��]w:	%�v'IؼG�iU��H�+(�Ó��j�=��-�,�X;��!H��9b���C�,��P4��޻,�H�H�:�Qz :ܯe��(�3k�Fa+�����#5��w�H�2�޲�߾�]���x�R� �8�n���l4e	#ۇ�!侩DaȾ�d��;�ɑ��p�JW��HQЇ�/3�Ǝ���;2�U�dl��8��Y6y�+;E;k��V�y]1d�$�F
$4 �^�?���d��t\���F-�N���!u`7���-���s/��c��d�$l�~g�Bf��K���=�[��.bo�P0;�y�.�&> �R���c�g�Փ��.��d��RVm��+ιah�xqa)��eR� <��R�t�?Xx/�VK�62�+�7S�?��.���@�h�ӊ���?��a����YJ�OG��2��(���%��p�u.��\�_��A盭f�����#��A�k�2�DxD}�CC>8�a��S@�w�E��ԮPEUVs������u�]t�� x2��' ��~���
�N�IBw5�z���g�$N���휻F�ةyI��P���[$Z�e�m���b��ORxl$��۸Җ����X*��׎��r�tK�l�I�"�э�!��LR��F����H�e��f+I�<��1L �/���	�`��&�3��:�M_�M5&�kkޓZK�#_Z--�#����c°�?�����9�ю���>��(
�H�W�9=� n�g1�E��	$���,�(8[[}��)��U�=�."M���o�ٺ~k�� ��>�����q���J�=3��d"�L�F�����X�i�2��?UN�EMx2,��V�i2f���~���f�t����T����e�B!��� Q\�2"�β|�9�qL��І'�Q��2V����,��,�s�ǍaUa@���5����`L_o��t�жM�d���}�L�)=�]:�*����wa���}���qW�i�8��cd��*+
�ze%� j3�r�/<�bSi�_��I�j�7J&<�bZ�%�ǻ�pF��(Y�����D~��Y�Q<��<�Tq�����9>\Eb���Q�М���Ţur�A��Q��g�����Wa�h����T�g��M�E�1�>L�@%����"��ٟ�T���Ͷy�+v���m{�	�j���Va���>BrT ��o�Q���z�����뒉���dߘx���>	����/�	����i.;xM�@֛by�Ϣ����us�����*��Z���tF��F9?J�-00�﵏��Ƅ~E�����{�ku��Kg��Ô���mi��w����(a��&��ƽu�:���z�
P�����n�饠D�&��(*l�`��{�L�(7f���K���?�l�^˿�3/@�}VY
_)������ǝ���C���
[�][����A���k��]��ϖ8���Oq�E��ӽ>D�B�QX���cd0�-)0HZ�����30����ݷ��PBj�0ʮ��l#��x#����|Fbݮ�n9�\������v��36�j���.��l�i��M�6b�M�.�}������}j�n�GH3(]T]m��"�p2���'!�I��vkj�o��Gh���>�Y%`�$�ZS������ALc�=���*�c�'�u�w]d�OX+�9�[r6[��̲y��ƫ��[�\���!�W��fld�t�a`���@3,��w ��4�9�������ap*8vLc�0��	�+mN�2�֕�}c}CZ�v����Y�$4��������3lw�����n�B�o�"r���1#Y�OܴE�C����9����l[2=	c�b;���l@�V(z�g |`�3s�T�P�����ԧ�A_������E��.8o\�b}j��~d�G �$�Y�C���j�����>�:�z|����=}Mmu8��Yk�NR*�aÛ����������jl�����!���C5޷�l)@��hY��I�Y��nΣ��t�u#����q���薡+��G�`�<T;k]:R�X:CNT/D��N�d�U'ԤM"��N)'�Ljp]Ry/ �=M0 ����Ӌe��Q����ߟ��e��W㋙`E㺃*�w�>�?�� ������$�%�Q�v�xZĊ��E���Թ�r(Y�0̃-8+�"��G�5�o�=�I4��b��3�],΂V�b3�[܍M�'�Fz��������n���;5���Dn\��q f�^~L��;��f�)��K/����غ7�
��`����.�q\�^w��f%��D�m�ޏ:�W�*9;�]@���x��@A�x���?�&9����0���5>I#���������_:]��S��a����u�V�3�Zf}Q3���Ss���R��Z��_�j�����)��#�׶��%�Svbԇ�Z0ʁ�Z=Ut�����lp�q��(;��-n]7!9��<]�E=��h��DY�$�nܭ�W-U��7*�D=���;u�R ��l�Zk�K��:j\8�o�����6K����G�6��_�b�#�N�k����0�f�d�>��J��ʐ��wn??Ov
��n�Mϗ�!�K�2^1�~&,��N��R� UL
�:�*LZ(E30���i��)��qZZ��:�:����c��Yn�2T�1�Uu�et�P��_
D�-0(,ܾ��QFz���ȋ�$��qR��2�3%s����(�^��u�P's����H�a���5���C��`�`&�����G�x���)!��|M�"v��^fvL�r�$�\%}SE�	E�O��q��j��0�y�^�skm�Σ�S�dU	�_h*{����A���|�w��ی)5d=�E�O�Q��$�`;R7�(�{ݖ�����m�Ң���k7qR�[� ,zI��[�Q*�N�`����g�2� UF���y<T�^�T6p\�]����y�z�ܰO�L�(K^��S����
� ���|f�"�s��I�L���g����CԛX�� SН͆2���Zh�X��x44�������
�G�W@�y_�K2�a��h���R;��� YP��� �q��'?�b``
����vy�)� B�dk#��>qX�q����7��<��W�2@<H��ސ�j�$XX�ss�x݆��c�a�M��n��}����Ζ�ߒT=��,��ia\q`����9�����+���*��XS+k���i���r8���� O�Pѭ��{�[�^�9��h��� �����^ӻ�}��N���t�w�0�i�'`�[oް	 m �$�34��_8������Ffs�i�����t.��5�r�r1f�~����B�=e{XJ�c݂א��B��=��}��t���8PC<7��ƭ��r�O�[Ÿ�0�϶^h��Ÿ��W���|����I�zr���5�01���d?kKs�I�6�Tc{�,^]�%�D[��䉳J�����B�y�6�\s�h��_��NR(�������U�����V��.C[uS�F�:��5���ǎku�UYKa9`qCи�'#�8lPe�=-I5�Xu!C�g��m)ԡ)��5XhE�HĘʛ�%���J_�re=Wj ���X��gNx�`����㜙&i#!C�z�/�bR��%�3ܷJ�C��Tw� �N�ݍ�Q)"���h�6�F.�{��]A�� ����b��٥��he�40+�[��y����Z4�9�����s�v|ܚ��9�G W�>z�����34UY�om�~��,�胚�<:�'_�M�K��Q�pl96��2$��N�
d��#)|�Բ@Fe��tQj-�����A[=(`&OF�aDd��t�	���w^oNL==��<n�p�]q����\]j�e�����K�R�3K\� `�o��W��y?��H>@��C9<[T;���ݲK�|�:4��K��N�T��U���s�Ԑ�[&��մrG��7��\Z��&�k�����\2R����h���A���q�$e򵠘��~��S��Z��1hqQ��3N6��H���}��t��`��%�R�ڥ�r9$M�*������ȟ�'G�f����!M�����I�X�����G�g��n�Kmo�2(|mw���xOLw�B�}'U��JD�w��Y�6�W5?$�n�g���W9+pI�:���y �dw]%v|�h[3���=3���f:F1�0h�pE�H����L�P7>�$a3��� Gx���q7��ꉏ�ӗ�,m�����||���J�˙��Y��g�-<`��j�]��b�_��t�O�����hZ1x}^b��{[B��%��#�u�b�i����gNn�c��JW�V�!,%���b_�I�ʙ�]���	�d~A�Ip�����7���M�����w0ڨE��2�;d�ܐ$�9d�>��R�k8��E��޸�;�㺄y����������Y8�l�����oaU��/|���x���'�Y�hN�HO�����J�Go�֫�����\{��e�ρ|I�($W_?�nT�:#'����W��!znrN7���hqC���a���}��,��Fy�f�x�bq�<.:��!����ݣ���^�`�q�>��"���`H��Ĥ�|��)�'ڵu�׬ǲMT�*&[Q%D�Ň^gm�R=���=�H�	����U�H��!���1l�Q�T0�	'"�_���=ط�%e�A�]�)ґµ�:�Q�yA��§�PmFלr��;�vL�t��*�飣�֏�Z@�^\��dЈ���M/��"��-/G;S�\��\�{yfQ���yD����ښ���$�� U%|gʰ:�!��ٓ�#��(R��ƍ�|����<���ނ�Pz8qb��SAk=���c3������>���#��
����p�-��\�@�~�{��@�~]�,(�ni�i�T[(��	��ӵy����%*JE ��^�G�b�%�����>�*׍e�u|�k��N
�w�DT<�id�r�&�p��C�m`��ȤK?��r���y��KM���|����$��>,V��/�ח����]W���V�8sS��gA#�������,P:�z�"ܲgp����������6윽��%���M�U����X��p�Yom�q�X����H3�3&V��__d�W����!V��{�n�_�5@P��	����]�[V���J8%���wB����&6�y��Bz	�\�DWL�(��܇��y�[b��מ�����R鞺�c��%Ҧ�ט�,�-��Q�,��U��mOG��h����Ʀ�I$�̎5=fm=���@�c�x&�EI��t�f��R	�v.�7V2nÄ��1��c��n9tD��_��{*2�̌9�.r�R㸍��W-��\a��
�7��SJ4���}TG��*�eEm�h"!J>}�;G���Q�0��g�KLV[�A���׉UN+e�b��v�@V7&y7Yc1�z�-=��I��F�Wdt��,��Q�	��o�&��U?)�����1�%�5u�F�r�䆴�����Eu��^�v�O
<7��T�ߦEQ�U6�ɉ�ܦ�{��M��-��!Rȉ)��癇��cn�`2z�@����\�WF:�����kN���>4�l��B�^o+]H�'����T��χJ�չnvF�fa��%�腃�m_ظ��(�_<�����0BT>sem��#��M�H�� �Q���|�o�hSڿ��B&S�E��zs�Ftꭲk��5�.˹�[�_ƕ%�\W�@�R�@.�xMZd�#�b��\��q�vU^��UA������r�.���cy���x;}�b�&�#�O[����V5s�j�C�&m��Ѣ�)�21�ml�M�Y�
�r^Л���=>�?�v��z��
"��s�Ȗ��e��]���Ю�q��?�^��|f�'�N���`�_�T6~���Y���<�����Ǘ�򬺍,�	�VHy��?�':f�Sb�K������P�`_j��y	o�y��6���.(�R3�<�	'��>�f�ִ��;]R<��fgr�3H����eV|�-��CGT�5��s�D˕��\$|�
�Z I����a�G���i�i�O��N"qݾ�F���D�ׁ:X�
o�ՖTE�6տR�̕[q�i�}� kf�;�Im�A���^͵���Vb���A���^��yO���Ѕ�M7ϜV��ɬ��_|;��ݓ^��@�:���_����E�ț�;{���N��9�fض-rڭv�z���x�D�T�����������Q/��~\��[��!R���_�By���vT/���l��#	h����h�J�\d��1!�b�L[c��+3���Y��~�BKx�&=W��m�����N�iZ[�C�D.y#�������_���u��?�y��r���Ӧ�͞%�.J����}�7!_�״��k���?���
_��5v���"��,(�wr*7�"���2yv�0t3WB� ���3��
^!�C�� �|w˂`�y����\�՗b:+�8[}��o��s]Иe�ſ�I�ϥ��m)���*�?���O�.�e����AT�Ju�����YM���� /��&�O����h��oi�����[Y��;��<J����	Q��1ƥ��C��F���NB��{��=���}ג��T@��� ���͸5˝y�vn��{��rP3_0��yI���v�0�lw���#%��p�U�]��+^L� �w�� �=��pEk�cd�5(�b��v�^���ፀR�gI�u2v�?�i=�1�P��(��_|�9��+�ݐ��c<�rp�Qo�Ū>�Τ�Q���7A��4%�>1br���������XG��A�پԒ�.%��Q㋦׳�r�5��f��x>.��Wy5�� ����xǗ
�CP�2�m��ÖÂ��8��8���Qo!u=nN�K�w���l�?G���]y��͉���K����������[Ƿ^w�FL�I��]����A�Y���wty�M<Q�##��r�g��Z9���*�̭H;�C��9�c7�.Tj)�ҿ��f��!4C�����KƏVu2�n��1W}��=����S���n�JԮ����0iOQ�2O7>��f�K	�=����2����$��W���
=LH�����49�����h�,XGl��~�]�JR��G��U�t\9u�b����}��{a+�Ͷ�3��c�}��W��8�D)�q#Bo�{qԀ�<����\4 ��6���O�1�=ܾp��I�6��:ahT�q�<t��h��QN-j���g�<�Ռ�>;!MyƦ�.�N��x��9���CC��U¬@Ug�b�N;�#F�����,��Oo�<��|�/H��`�L�y��8��	7��r������q�(�7��#aB��yg��,ԑ;�)\U��S#��E�<��1:�rP_
�7��*DX��03Z$S�0���a�@S�D���"8�'3���ֶ1�
�UX�`���.9[�A���:8�i) �7weӾ:���lB��r�{�l�o�c�d�$�ߖ�]���2�K�*`%y��#h�6�G�z��%Y�LPԶ.Ն��<~�y\��C���]/�1"��H� �H�S�<m�R�g*7����r7|N<ѣܖ /d�W�=�Uu{�|�&����pG���_Tw�4�Nz<��,�a[xxd���ʦB\��N}4W�`���,R�b�~ί�83������)G�{Z��!U� ��#����4��c�� ����7��r���K]� `�� ���/gR���ϩ�bݸA@:�D���s}kl$W����\��W_%��r�*|	hh? ��7T��d$��VC�,�4~�~t�z�j��q�n�F�}��6�o�A�"��<4٨\���!S����s�TGC��rʙl�lU�u����b�@����}ec��H�B̜��t�}s?fQYvS�v�Un�"U���/���e�����եf.+l6	�.	�����h��!�4�8!�3hYN˾�q.�>e����(b��B�8y�и���*�3����seτ�6|.��4��+��֪�73��'[�"��^C�ٮa�1�v3�}��/�Վ����%��&+�|�"/$�E	<�7䋺��q�<�/���)�zU�N��A�X:���xŷ��!e��V�DG������0&ogQ���Y��M����O�] ����O����4h��A�kF<��ɷ����;ȍ;��3>(�O�PĂ��[��ɠV���&$��b���r�����1��eNȉR��f��1�<蒠K5g
D�]Ԋ]��&�N��谿j���3�z�ȝ��E<��1�$�G&��K<G�-��	Ac�$� �7�M��r|�R+ü>q��J����0��FB��g����]�W�Us����-'	�~�L�y}�8N�:e���ͧ`#�u`X Q-�C���5PM��I�Q�6���{�B kM�Όo�U%���a������Qe�����>�lX3�j]���y;�����`-Y�
����|`q.Sg��&���-s�5˓0����$A�s,�� t;ɜ���̳�4���/eFB���!�� w�_p�hU$�E�"z�K���4ׁ�k�J�aCd��/���D "�%w?+4���0��Q�����w��:I�-�60HFXy�j�;��S3�'ĿQ�i�d��A�	��U�o/�U�l\�����3b �@�
�38�]�Ju�A�/�XB�_�D���{����amA�@��'ޓ�R�B^�����	H����LI<�䪔��I�!���Ꮓ�5VXA��Ar�[s�f������C���P�AW�w��M������`/��sm�q�}���Z���=U6��o#��Թ�� =)|� ��P0Qi��NP��rU�š!�s���¸w?c� $�tf�!��'Ց��(jе�ٸ���D�F��q� �����T+aY!�uZ�c����ߌ���k[6�'1	t���MOQ)�l����+j�|9X�M�v�^�D��]c߾�&�W��<�ܮ�袝f����Df��]�ƒ��k4��>��7-e�)� i�p�:W@@��瀞	��5�s'2��u�|���(�i�4C�n�F��qv����XF}TO1������!�	�ݷ��M�E�A3NZ}L�BO@�C���E|���L	b��kO�򱽅����86
љY&ea�v�DoBe��;]lg�!��>�+���� 8B��tLB�(m��Eb�*q�-�7���w�@��B��q��B�3�ܬ��ڂ+�Q��1??u��KHb��wן�E��{���A�U,�4�~gZ}���8�
����ͧ��Sg���m�6pDJƦf�A[,ʏ7������-�(Ey�Υ��	��ʓ���f�T��-�#�NF8y]���oM����6��.y������؃H`��]�'FNKa$CMr�l�j2�1�D�!��ju<Xz	?rh����G}d�HSm�MK�IuܠE�9)�i���x�k�5QM1^��2�a��F�����ə��8�3�.�H�J&U��Z��$fn#W�* ��<���C������,=�E�$S��A�Ց��v۱>���L��'�I���u��||�ue����-���'�1���G;����.p���R���<�.m���^p@T����D��g$hʏ_��e:���"#��X��x��m�ժ�w�X!:���Ě̸ԶP&���&���hVk���m4]9}�� �csq�f+^��U���zu�?FGp��x�T]��F�HaT���.t|��.(�1���%�R��g� 9R+}ߴ�F��CT��:��5��3t����r9l1��^m�許g�������3���J<�E{�C�D|�d�y�N��F̲o�4��@�@��vT- ��@��']�1ĕ���N@ueg/���Pa�~P�Rmq��a��&�O�[	��-+���,|���ѻ�[n�~�ؿɘ���Q��w��j`��+��b�qS`ұ���h�J�W�<Q?{ؚ���VdU��7F�R�Ux�
���C��uB4�-�[׀���W��KN��*�O���o��{�k�lYx�|��Eb�ԛ8�􍈠%hÚ��Wwox����}��(��Ƈ�B ��CK����W�¶��@�d������'bB{���c�QN��g��]S��d�D"�ޘǰدgx��u7�<�Q��E|ػ�p7[hL��r[C��5pW�� $����~]x4;z)��#U�z�E�w �\�s?%���C]N��
B�Z�V��h�w�CY�z>�/�[]1Pe���Gf˸�s���e%]k�w�T�f�:4��ؾ�jT�ܩ#-H!�H
]��D�V_�%�<�,�#����F�ٓ29�P�m҈_���!� Z�7��Ǹ�%��5���a���İR��M���/���>�N�j�2�C���ٯ8PLM�������	](L�^PR;�Iw�`���Y��P	Kw��Sn rG{�j?��D����\�E#��2���h^QJ�S��C굣�2iD��m����2"��ze�v>���|�|(��o=Zq^��n�v�-ش+x�Fc�u�k+����s���]<W���9����Kz�7s�p :�yl�|�7h��5��p�V6��i$#�iS�a�An��L�^U���l�^-�V����O\�G�~uQ^���#ހe�i�|[ �������o3�U:U�㙧�c�D�?ϓo�����Es#S�!�}�gv$�/���i�${�E	v{��?Q�>���v!}�M?���7��aP�Lat�4`��B5©y��D�e��<p$�	$kI9LdGs����k�`�f�w�}�WO9e����Պ�"A��Y4����9��?K�+9Dc7v��ȶ��] ��	����m��	�&]�ІN�d4Y�~���F�Z�x�� d�����\V�0'�<l�� ��\�D�{&a��NY�;IU(,ڊ�
WpZY92W��&g��/���Z0�,Ь��Y"�C� ��UP¥�' {|�Xk�.�E�I�z�â�np��4�6�)˺�U�EB��e��J$P�/W8duª�m(`=�H%�˦�u���A���g�SgB]v���9g]Z0��O=�LT�6���v��1���%��~��D����Z����������}~v�UB��=Z�z�~����>�\�jh�N�5u��x���cΨ��r�`_iϗ����JN�(ޯ��҂�Lw݃�t֧��j���J��L���Y��>W���wn���g��mC:��w�a	ßM��)m�%��:�Ր�Z�0��>���X��������L5`����leF)���-���B(�t57�&�9o�Nih�/��u�d'��3�k[Nn��C3�b��C��M�g� ��ॸ�:xh�`��=z�Cb�v�&��s �i]�����{�V劌�9���X*� K3��3^�����LHȊ�;R:��b1g�ꢭ���g������`�������j�Xj~v+���g\��Pрz�|-�|�* �ԛ�y�˩�9�/�[�_�鶱�6�W���.#�Db�R+j���h/��J��F4ߺͣ��4\�[�% z�<&V�jiL��q�Ll
�Sq���}��)����>k�h9P�!���.��(}�����M�������9�d����5��w��$8�c"���q�VA^�{���g��ʊqQ�ʖ�)M� ����"�JFᙈ�?x����4W�����1 �g���i���w�W\�.�c���rIus
_�~�����?lL�����A��� ��J�:!��	����;��,0�M%�K%lL��}��������.=��"T���]k�H�2�,N�'���8|��ˮ�t���lz��<���G�c���m�%��0K7_���r^&���D�ճ�Ti*f����݇3XU��1U���CvdN�n�����E�?M)4^�F�z/�y�z6���}cVZ^�ϼ�)�q���`d��������F?Z��sj��k^�©GxߗB�@���8����ib�ۅYy�hJ7x%�3��W�k��t�Xٗ,�7i,����0�5t�u3�3҂4(���,�m��f����(YUIy�p�,����lP��u��e }����7᪳H�+�5)��4�l��k��ǒ���a.\<-�Їh.�mA��TS����>T ݤ1�1�*����ӑ˵9�0�)�}H��_�ͬ�#�"�`%�AnK����:]F_/�ѻ�N1[�4'9(�5��hδ���MA�2|�6��-���V���ѓ� mm�,�dP�Nc����U�����@o��t�
�p;fu��5�-޴t��]Lm�% ��\һe�m�H��E;�P�B�Z�s�)C�^��naz�y���n-��O�����D�'ِ4�������$Y�=����
��#Ր�@�iE���6��%%���^��Q������l����uDZ����l/��`1Q���<�C!�+�e��Q>��V3[�A�y8H#����_�|�MIiFc�-�%���!3�)zS���nV��[�\�(=u�m���KU����9���J��:��{8Ŋ�����Θ���-��kV��D��=�o���h	j�V�ih�B��PZ�`��K)}�̍��\9T�	��2n��$�����҃�6���\��&.ф4q��=�1ӱ�����w�_N�{i�8���{=:7���w;D������gEד�EF-�'u3�@�3c��1�ĸ�E��G��m2��"0��F�{���];Y��� )+}�Ҕ��8�>���<b����26�\d�c����E�ț�K�rB�t9�r�B4�� 5�A�yӺ�Z�v�w�@G+�?+UxG� �yR��A�*��>�a�pP�n�B�`�.e�ɛ-�J,9s�߿�7�QJ�Yρ��n�ց9�T�d�Kr|΍��q�<<}��i�r�R+=���|2���N����0S����:m}�2W��U�z�Y�s	�+�,�S!�]�F�� G%�+��3�h�����$�wΦ�V��-�R`�g�������IUԹ ̶�J�O�o���+M�fU�A-���*d
e��N_6��>@�f�羨�z�"O��͙k�+ѓ�F>h��!���� ��������N��;��m�I�1��h��px*0�޷8'�9�T�ȑeE�*G#Tq�]�"��}w����a%��#���D��_1�=���$�f)�)`��k>.υ�t������KWgy�s�ډŮ��3�N7�8�p��YηƜ�x�V��QX��������#c@M�$_�I��>@����gqo/Y <�Cݻ!�^�� �.���ڻ���vc*`@8aGO�s��l�/��������~#��a����X����:����Y^�K�*8����=��e��1�#�O�@�	���m�_!�#�
X�qftȆ��^�*`5�=x�~���e����Ѳ���"��vueK��e�
4�˜�����X26�\%qb�v�L������KsZ��-1~���?F���.d�G�� y�(����^5���K��������< M3tĮ+Bp��ե���t���?�Jd�m��K�P��2�XY�.��q�~F"��N�h!�X"���c�ۜ��o@�z���_�0Kd�d5e���qح�S� ������R(�y��I�T�����ˋ�~#�U��n��̲N���� ����?�G��W������e���9��R�Vx��F�����>�Õ[�F5�^�TI�D�4F�2����{�k�Q��:�e�Ur?S�@9�A�J{�]U��߰<���B��a��RAX'8�.%/~i�5!����k���p�^.���d�$_D�s�5 k����VfZ��<��z����>>�.~J�}�X79H�����n�n��ј��>�}������������o���I"���p�7��a�l)<z�j�q�6��/�Jp?H�-��&�>3~щ���~\���b��t�;Z,�{���.���#[ߛ�Zu�~\	�й�L�l~PM�܉�O2��-!kz�ǩ����.t5�1#-�HM��X��Q妱>����Mn���T��/��(4J�Kԧ�/�#�hxI�<bb�Yd4)ΔG���� TivS����tn�#�:X�;BS]ЁJ��Ro�0zU�]]%zy��ծ2N��P�M��O��zb���2y�I�C3�GС
|����<ê'�tQ+�.���Ԟ��4�6�L#8�=v݄k��Q�Fm�"g9{d�$��7X͟�&:��g��8lY���%�z*�/"�p��I=�U����z�묐���b�}Nr	!�o�G�z��E.K�X,zd:^���(5pTŔz*g�uH�{gX�>�p�Yh��Mo�)F�T|Hl}�M렿��F�H��Z:������{9�K~G��DN� ��}�+�+�qv��8�ۤ>xk�w�\��~$�jQ�~���^[N���� )ߡ�CZv�?w7�j�D��Qy-�A�W�I���,Jǯ,�5jO`Ĭ�6ZY`�oP��*�a����9��Q�"}��J''������űu��{?��������I/uM�4c�{��������Ik�ߣ��fų\��]���+`_FYq����Ρ�R��
�`��*jl��n�ޡ��T�T!  ��7j�N��e���F�Ѯ��S=RC��q�҅�D���[�Kr:DR��~)�F��)U/y%7��ju-@�<����#�!����-�v
;#�1ES��Z�D0+}�7%��^i����C��'��C
����.7�O\��60���S���s��Y�\����qx�����s��\�X��0�C��3�NO��:��ɐ���Tj�������{J�5�EW*�"J��o:(fХ��&�Z�ǽb�Ao�P��m��G�Hb�9C_AI�rU��MK�#��d䫶ЈB�`�	�'�?�^��~�tR�>o��Eږ?���I*���uӅ�}�������z�@���N�5���#*��AP"n$�s�&hp�V��̟����u�����q���!;�:`�$A3N�[��5_l끒"n��9�g���ׅ u��'��WC�T<��H����z}=����W�],By����Ȅ��3��Jj\��@	��}������g@n�L�x%;XA������A��ATlV��+��F+p8����w֞�yT�*7L[�11��6���gղ�b�>Xɶ��E����5$���/w������������\��R8a��ɐtcxx�H�As 
�q���V�u8vr�41Ɯ`|+2|��">�T�줕��,�*[����)��-�2�t�����b<E�#B�˻�+��D��`��A����X�+�)S��i���Lb*
��˩�>�1��)Z�i
.��N`K�=젅��q�yc��	_�G��@`\^�:8�/��S�,���K�_�6S�I�(�@�h��Y��,{�N؁d�!���`��4B�5�]�lcl�\K��>��j,c.ɻ(��(�Z�r��	!Qh�}O�HkM�@�2$/�\S�4��`�d��wz�r��b<NbO��'�]p]�m�xui��be�}���w�>�ϵ��n���w9�.�qb���WMq�����B'�LJ|_���Zݛ���@�0�9��|@�Nϓox�������>�1ߗm*��c4S���k�\ �
s��ܥ�"��˦��C1�3�	L�//*�i(H�������JY(48=S÷����������fE9/��.��3�Cگm�n�gU!�ߢyt	��p�e�,��zϻ���暊��e�p���.|!���7"lz��/;�[�`�O�TVX��=�e�ڎ��	��y���t�s(9���sB%k0
M�I�Tλ�1!�G�*'�m�� ^�"��ˍ�'(��1|�]`	���L�Z�i3��`Z�q;L���Wn��mA6K�e����V�W;K)O�?�I~�nVNK��\K����M��v�L��o������)*��?F#�S�A�f�%�΋�7���ܗ�O��U�Ą�8�9��n�[��n� �۹��BV��ƾ��(Ԁi�y�]����N.a�$ס�mdE�{����>Mf��|cz���nK������s�ٷg��f�k����۝�p��$-T�6
��<O�J���Qq
d�5:���I�&�Fs2ok�$�8���M� EV���[���>��oHǫ�`
�k�[��9=*��a�*�">��UXa��u8�c���Ɇ�v�fV�����p�&�(8�����F��0h�:^!���Ҡ ,�!�d5��4[�JZ�v�V������P�;�������1��I/T$��|ľ#_�l��Z���Ƚ�(L����ʴ+��,E���('*�pE&;2�;�@ԭ�A�e��d�F7r�����}��4����|U�����'�M�j�f�Dk��O��~�	���;ET����8�"FH6�?���"R�B�>��G޷'U����I^�pI蠙m��=�8�(fT#w0,����^&R^�>B:c�('/'��?ǳ$��ٽ��<��%dH��di�{�x�kk%u_!_:��8�w�K��V�ͷ�eU(��.&�1�<�$+-��u�/��V8#"���.��`	��mu��6�ui����|�b�4Yώ�M�yڍ/tl/�K�\������9���љ�$M�cwjWXD-��ȭ,�i9�����`c��t8t��XĔ��DfT��w��217U�}�*z.U�e	6`���xk@B���hS[��l.U��gA�O���O���c�^(sfW/��F1=�nn��=3sx T�N<z׊�#��z'�ѽ�c�:�]�g�!ǿp�I������'ç���U�G�x b ��u#���X(oK½���88����̴
#��� ����uϢI� ��}t�(J [�P	�P+'?�ӷ��f?�}� jr-�𤈺�20A���/ �'�*O���N'��R|bJf��E��GK$>l��)��qQw1\�W�y��;�t|����3*!����*%.�_��7����\��ELz�l�3HI��:<�D�����*s��ղ8�:YB�>�A�<4�$!9	��(�G���RX�x�Ք�l!���)�L�J�K���`7V��gO�4����žt-�fm~2R|# ��.���p��W�R�Q�MJV�rAM3����viᕾ�ߣ4�����ܚ��]&��� �\��Ǧby�ؚ�%�©T;EhZX���מW�z8�7s��qOx���u�Ĝm�#�umɻ^�TMkJ�)�W��js�:~q:Z=J�=3���Z��LhNB�fo&I�#H�.m��=ϯ�)��)S������7��o�TRM"<��t���@R�w�
��ƈ��"��[�H��!pm��b/�=��D�I��V�!;���)K��Q��t�jE%Z�`w�U-�=��I�p��:���*�0����b�Θgi�_���9.���?��o��'x�`吐	�h1�̌LS����1�x��9r���C�ֶ������^;�;6>�b�v�R��{�뎳���9�.�q��2�Jx�b0�/(rd��5[Uc�&�ت�i1�k`ݜo� �N$��#��'���� ��e���V6�)����D�#Z\J:b�]�(��T����Wΐ���'���_������z�{�_�����q7� �[�q᮸�5L�[��#�����#T-��r�F_�$P�x�]�l���H�hI����6�Ũ�S�ȩOI� )#Ql�c�au���g�p&�O�<��X�]tGm�Y[a}3�/�:gG�ݢL�m��9�z�	w넪�@� �Vj4�k+� �������:�Z��r!iC�������4��dl��ݎ�Bp��G`1��C�g�S��Shl�u�3�f��u����Q�f#e֣;�.cG��$�ܬ���b:L)�8�����8��C�*?�Q�Pw!�\��6�ᒁ�.ࡅ��|T��9����ѠmPx'�9N&?p.�`���|�\"^��A�9m���~V7oB��f�'ޤj��x��=K�>�b���ѯx&�e�W��0�T1-��qS�	`�V�Jg�\D�� U��e��8"�k��l=d2��9�4�|N�c�����N�ZY~���ˋz@�'�%b1Ky��L�R% L.Φ�����������uќ�����+�tǽ�=�3����WUY��j�h��|�#�4;[0�z�MŽ�g�y��P�dq�A��)�K�r�o����H�����Z�n��i�Z�tk�]H=ٞ�\n+��OY� E����K%�/��)��X^8��Wq��(�ۯ����4��~:�.���������`]A����Y�x�v���(4��l�FB�AĜ1ګTP��ܗ�7"N��Q��z���)��뵗��![�qi�o.���<�BLd�j��d�%6�,"H���զ"8����W0C8��:������`<���Z$�w�[͗�������Ugh�0�8DBOfۨk����5��b�J'®�~�r����<=n���%�
��=ZB.O�f�QpT���� ��YW{'}0~Q�ݜ��<,�-�Ì]�]�\nv;���w�Fl���rm<���>/�P£���'$x�6���y��w�X����*Ro�g� ��;��?D��^�;��q8�]�ϣ�v���$$�w8�n�ϻ�C����_�lU���\)��S H�1�˺q'����`/�;n��DϜv�����L�=G$�.L�[��IE����e�ȥ		�"���т��Y�D-��h�)���(��v0� s��jc�?-Lxo�j;ȧ$K�L����9�x��ż� V������*� s�K��/�S#k=��_E�'�I���'�
�#;�i�
�%)ߚ����gh�y=zp�"# ��lٕ���+:*�i��$`"J��v?�(� Z��OE[;��溍j.�fjUv�g�z�'��� ���65��f��~�~o��2Ra3�}/Yt��(8h��o-��<@Yl;��D��ޛaf��g�M�X���뺝��X���M�'��Je�w�5`ĝ�U����Y�bG�(���R E�+�W��F��>�FQI��1�){&v�I(U��2�����Dh��DH]���G��s� �Ԓ"�p,��c�D���^����Eє� Z�D�i,�Y��K�D<m>�� ]������C��Hg㑷u*���v�J�S8,28P�C�������8?�W<p�p2��qy����������O	�b�Y�j�0��z�+�>��֞)1BSC����
:�8a��}.�aOT�=�7n�_@�i�M�lҐ����cv��B������ɝ<D��ލ��5��f��4��Mw�x�2[B�,�.D�����˞Eaa�}��s&R�N[��l���L��������C8\ȼ#?rn��V�&�#)�uWR
V<��g�
V���R*�i�x��|�w�r%3o�Jc���4�V+[5����;2�2�NM�B���<{a���d���>#C���%�6{���K6�V:Պ�HJ���.���� �^���Fm�J�3�A�~M�9XusH��2fBM;��Q��w&O�����c�D�C�g�Qi�J&�.����L:����8�rU�\�?|(�@Z���b@h��g@�����N�sdy^㗜�����,�P�8�֛��Q�ȼANT�|dh
�E���8�Qv��G�o�cG�}Kߕ�[l]}�Z
fw�#8Mɟv�Nj�Gi���W���]�J5��] a.�cA�����?����<UQ"tߏZ₨!������n��ԏ�lp
�9���/�8�p[���'6����4�ޤ��/n6]ͩ�}u�w6ݫ#�o��YC���p��E����]�X��H�B��O��t-����KX�Uհ:w���I�&��x�-
��r�ņ:j�]ո��d���������e#}Jt����Aܳ�m��L]]��@�~�,M��cS/�ͯ�<�ٴs����*H��a�F7e_��l�u�iU������w
��^��#���\�U�5�"|�BN#���AiA���5�+(F>(�L�Sl>s��WP4�^�Sƶ�<��GX��dړ�,"�gz�w�8D�`?+瞞â�hBK��?4���	ྭb`��'<%�+�̂�����<�D��L%�w�VS{���xV�åVNEjxII��X3��b�?�J�Bo�|L���Y�/-񋮆T[�T��0%��h�!��,���mn8���j�H݇\l-�Hډ��BN�B���ks�gi��"�����w�a[.���ݭ���׉fO*�H�U�4.}\�^�m~���5.8;%��� �=�=��"��y|�BW.Y�h��,��T�'ILd�(�̅�c7���t���0��v6�RʌG�#�Q+�=f A��G�!?�=�"[R��l��ZA�� ���7�ڋ�d��Q�_?*����޸uU�אM;h@>)�x��p�8��v�Բ����Z��/���ƶ3�ɂRokA��,�?!�ƶ�̊+V h��с�@.e1�u6Z9n�sz�T�b��~D�)$����!���9����R�,�9=uUN�>�zM��}g�IG+�>8P�,���K�PW܀�Xڮ���X�G7w���Hm��e��I��|����o,�zk萂?�&q����)��%S1�o=�)ో$ ΫX3;�+K���	�\�"N��	��z�Pm6���(i7w����
6����3�֔ M��pe=v�6� 0�`�M��0�������ãJW5�[�a^�o���)�jȴ}ʈt-�y�.�|W�-�)]�n=Eqwd�wo���'��3�z��B~�8�)�u���L?Q��}��}�6}aO9u${i6�H֚� �vN�D?���C�`��	w{@�6��̯�~�v2��זS����b���a�r�@/�s�H�=*v8��H���C�}���:�ݕ���֦;���zd�ڑS������-��n��Ƥ�P��A�*�EF�
�����ftL¿|�r�y���I�4��1]c>���_�#�Px��� L�qF��%ZJ�aɇ7џc~�5k�Ǩ�
3��ƙ-��;�G�| `9�"틗���҅f�,��GS��8]��߭�xd���md�;E<Cs�"�����8;W[��p&;c�����7�#.���C�x,�w�IC$����u0߾\�<Y��|��놐������پ�*�&|�K-{�>M�:B{��9zʱ��k{��l�ғ�� ��+���7i@�|E;p�!6�o��?��^�'|���>�cMM�[g諸% ^sc��\n�X8&�@ �jt
��6�i
͖"T-G�6��n���C$�䪨�#��ɳ��,*=��������#,��q@��n�"�"�p��ߤ�`&���E�ݭ��c5M7:[fH��h�+��N��@���)�XOg�3/.�<��Q���e���(����8⦝�l(X�	o�M#�}uiӵݍ���$�tY�-������U?�3�l ���E�L��4��R9d������=��� �P�2�I�k��_Ҡ���^�}_�B�U��S���ki�z1{}/�&�$;��N�������^+����k�
�L
K� 3���t��oL��6��WEk4~��JDK�xq��:j����C�!�ͯ���x����������ὩCҸeEuW�Z�+c+�{�m� �4�y�ѹ�`h�p)b�
�#*- �m���_BO�K������~1b9����s��[�Vshͥ�QC_�V�v�_v"A�o/�CL��ݟ��&ֻ�?!�\�X�i`�1s˿��[׵D.�7�j%Sr����Q������og�FqL�	��\�|�������ȧ-�IG���W,(x.-t6>� �V� w`���C�~�g/��B'= v�E���n^�I��C���������+Q�lR^;S><b �
ZJIwQW~�nv��|T1Y�� ����c�{r�KN�Ы�J��	r	�d�pm��J�&E���`�OJ�<����4㎓�Tw���A�vSiy؅�)|��L�c�0_;z�H���|�E�^Sz|�����*�˫��A!���j �G��9Ý�:(6t ��$2��.���YJ�k3��꽚;���2���6��^��ZfL�g=`N�8'1q!�栌�hEv8AAl`�kK�QY&c�NU(z�jj�G�HX��ow��"�&���͍vV�`�J�wD�QPp��"϶�w�����tc$��PS�����]�owI�_������F�bΆ���q[3�g�Hi6�$�V�ں�ٍD�Pu_�����<|���3�9��	.5j~���Z�b#�q� �&
�9!�v��1�}�si�v��ѱ����E<�
?Zsl%D����t:|��9��1��(�Up��(,3�P*��Cm��џ.�\�<b�ь��SZd`��I^qLO����c���7nyQ@��s](��R�|y�Dq4�-ZD�z��:��؎��[5�J[G���H�!~�oi�f� :�yN��M��|�����/DQ^n ��awh/_���J,1!�#<�f��$�K��UK�4��Ȓ�&TK��ef���]χ�]�̡k�Q���F�k��^:S`hi)�����y�u8Z��g��!�AǪs��j�O:�3I��ˌ���;7j��^)n�`��-�6	o��a�^������7w��:�A�p���bT9�e"�dݒ��MMx}}�N�`�A�#����J	�k���/��r�D*+7"�lE	���oO^��ʬ�)�ӌh`w������g]@��"+�?��jQRE|��&��d��n�%/ƶ���D1J�\@U���<� �Pq�7�U�*�Y-�Й���f5�rzB �>�ݰ����9/��
vg�@��a2v�;@i4���ɠ�C�q�y�����l䨱�D�M))�0��A6r�k�٤5�u� �#$��L
k7چ�in��3�&�� �}V�~�r�Ҩ\�Z���k\��q���pD"ǯ'�����\+�t;�]�:jC^q�����m*�_�"k~�LY!��k� 2B�8�R��/҇�8/R�>�X|�.� �u���'��.F��35u��X�!�4�~���� Zҥd�����mHF/���ۇ�+L���mjR�{�>ڈ�a�i����[R���N�?�2��r/n~���&��њ�H��v֕X�I�ס3�j4�[�6��pKu̡�oi�J�Z��gҹ���JoJ6F��z�=��+�#@��f���hY����}Tf:�NT(Q�m��q�i����}ˍ'>���U�"\�lכ~�F�����?�������*��zC�/~�oaHi�6*���d�A\��[��P�{�����_u\�dDϞ�^��o��q~+T����ʠu�/?�T�^Z�j�aI��Y���5<}��`�1vNqV��L���=�ͭ��NE��VT�G:��f��m@��9º�hkn��HI�����������*��C���(��(�c���"��z>-�ѷ���ñtK֙�dc�+�Ӂ�q6�=o�����S�H�u�����R�nN؈�*���x��K(� �G�OC�`׼P+�]��G�P}�7o�K< _�ِ�iZ��P	XD;���sI�z�}� /���NtKT=���a^�0�T�A����"-%[���֨�_�J��(�̵ZE��}D4.���I�����2�Ц�)��k��BU��6�
!�	S`^(�E'�!xA_�V��l�k�S���M2�>��W|�g�F�EX��,m����7�Fz�E�t���"sH;)r,Ge���&���뼉�N�FoҌt;׉J�b"���`6Uڡ[��Ŏ �wN`Q�D�4��e�Y!���wE[�va����XJE����P����ZP5ɊH~�aI�_�?1Qm�gPQD�09�(C�F϶w�^{�Fpl�8���:�9�r�Nw�����:PZ���h������֒��b�����*׭�3Ը�u�a� ���k�~^��|t�w|вZ�+�t��������?���moǀ�GZ��^Е�*���ژV�D���ó{(����]�t4�=��0K]H�fcN�dJ
_m(1e��ˇyv��`'s�v�dAw�XA�$ �e��f&,�9�{�Ҍ~�}����]	�Be�k�R8@4��e���|p�ُf�+.����F�K��0hKѦ!Mm*w�������\�R�싵��	W�+W��UR'o���[[B���2w��|���+g
F7�aR��zE���Y�"wP�?���YD�5�t�/P�%��s;�@����,�#N���P ԉj�`ň�\p:��mpicGX�{^���KN��,�J+b��~d��egT%�uG�.�	V(�������/��Z�p!,4���n�}�,��C#=�񷳦�4y�������c��0��H6�)0'�J_��us��9p����Xa(�.zr��ż9-(CI�.����^��;k�դ�~�Oxi������P j�l!�I������M5wA)��i�x�����2�/i�(����R�SS��9TM3�R��*x���ѓk�Z��J�?�c&ٴ��ZTԫ/�ȵ�H-��s�;�Ӂ�;�U|G0�A4�T%Û���҂_�����8�{�3��4"��l�+dKc��o).�MmY sڴu1���!�5*���Q�[V�2�I&�4:��懂	g���u#�KW�m�$����Ut:FE��wC��c�Ve�U�|���w�jGsy:�+Ĝ�*�}B8F0�# }8����Q��n9��➾��W����[9�⡕
�î�:y���Vt.Rѐ��N[����-��W��x ��=�|J�"'P���ss$���;,/ٝ�T�u{�Z�QS�ML�v�W=a{v�b旵�>3J� �Sg	���ܩ���2'��]��].�OL�>��nn��ӳK��f��q|N�%�c$��(�t9}�}�R�lwc��>�)�a�d�%�Ķ�&�K����_]�"ͻxꤺ��QĝF�p�*&�)��0�"Dӕ*��U�j�][�I�W��o�!p��ڭ�q���zTD�lSb��/�}��q�ŊR,��]g�8d�N?�E�l���XJ�ty�bWk���F�El���h/ջL�t�k���@n�"��z����Q5���F��=�0�B�-ɤB[�Jf�I���2럨)=����~@ �����Ɲشdy���Vz:�
�V�X��|���}mkaE����n@�D�~�-�_�`�;2��H*��z�Z�����Lt �3O֯zH��	dm��^����"N}]+���Y�ͣ�H��Ge�?\m����'
g#����U��bmXu;��Q�.s��:y� (�t��Gw�0mQ�ڔ.jY���{W X歲Oݶ�0�m�̧Ⱦ/7���&�2{PDy��f�=�p$��%��P�P|�����X���)���h�9W�l����~�Կ��vs�����d�N&��K�A�-�ׯ0 ��l�"G��:x̬"mfO
2�ڼf��8�6����7�)�o���&�����>c�^�N�Z�FEw
}�G䥣�s�	��~�c���|ri�PтU~,E">Ȱ�o��),�5��i�2
K�^��$ �-�$u�$siY�V"-�j1wݽ��r�N/0mS��l3�z��խ�L�&�n��ا�VPa�(�2�.N#�yٮ��<����d�F�@p����M;'@?:�Ey��۔�hiD��h����V�c���Ow��eVR�~s�L�9���ʧ����4�����Ss�^��q�Lǫb.C㊠`��C��#�K�����$(�l� �B���_	n3Ã<���F�j�$� W�J��=/�/�a���f�w�uJ���Y�K%�xc���EAav ��փ�>��wx|<��"h��d�WX_�_@�1 i�/~=�<���7�������/�А��w���'���u�"��l�v�.�,�0`��J |�����<�p-�)V�ޕO1jh����>xn�3r��S��um����0�C'�G/���zS�� s�2��f��o�����qS\�����QW- �tҫ�ꁝ�Z�j��'�`�[�Z�Ò�N���v}LS���{�Z�Iqbڕ��=��QJ��W]}%�M�K� E|��Y�5�����/�f��؇]��qIS��;[+�,�������WOн�v�9�k7RG���$����v�+h�oz�D����Θ��We/��6
ۜle_�;�����A�X�'18�-�|����t�0��ݮ�^��GsC���y�L[��^�P��r����]�`�w>��ʶY�#O��dk��Ӿ�09�K�WV�Q����!9�nm�V�
�e��`��K��3i>������d·w⢰p`���ʾ�2y�6�
j�z�L��u�Wh�n�^���A�X�J+�ܐ�N�ؙ�aSv���텒1f�g��K��d�����Ыb(�x��c�_Dc]�j�U��oL���M��lQ4��="O�g��ٕ�����r��B�g�3�8̀��%x��Th,������Z�|.�)��Ȗ�d�0HHzY���!����^/�a`?�����g(�@�D;�&�w� -����e p�*`N���C7�dm+�Z�[B�֟�毊x�H��.� ʫ��S�&kKh'���QQ��C/��"^+=�:c�"�:�f+�`�d��ț�}��n�� �$�~-T�L�1�����w�rɎB�3 ����ld��M���l��H�/^���n��i�C�=��O��ќ@�^Y	���o�Ҁ#yݙ̀��3�	��>ICД$H5'���˂�L@���?����QC��ڥ�>Q��i��3���H���e����ZFJ�汣\�W��H�Cq�B#W:3��[��n��F}G�*(��q�r]���0��E1���1nŇ���f�?��f��H�1�`��.�5%	UZ�b�˖��~T�a<a�T1a�:ӝ߶!� i�e�.�;������=`~�����yD�϶x�C�j>�;��1������_�g}W-���0��$��9	���^��q"ۘ�$nK';��u���Ph'DH��s�}�������.A�V�ǻB�m�D�a��{,����:��T)�r} �+�.v�h4�"���)�/S�������HmDh✹���BZQJ`zFq�6�7�'|]w]S�:��Y���[Jߖ��o�7����`�n�1k&�(ŷx'�V�w�2W���qQ@_v`��R���!���ݦ��a���Wl&��΁�E�f����eN�g=�&z��䚢=Z>tR�g-k�8�xHn�/���w�!��y�v��TF���Xy8�����^�Q���HJ�S�e�$��t��+�_�ƨ�a��+���.*���R�A޳�{B�w ����iX3��k�)+I�<=���(%l��Q!{z�u���`iN��D�Lri(WNO.�{p}���_k�1+��l��N�H�4t���x�D�l�(�$�K��ed�
_9�M�}���{BtV'Nt�d7T`L��3�`FV���q�F=6�S3ʫ[ UW��VTv1gF���8�V���B=}��������Pdb(�9�И\��)�Oi����&��%�.����Z�Y�V}^~{]�?;��S�7Гq�+R��Tr��p��~m�j�ӈ���qxXɮ�s��_{	_1�l�z|��G,������~/����YV�u�[Hܼ4Gh=�!عh�D�9�h�
b�W�����a��,��g���RL��T1�&�ãl�
�e��
�0L����4�s��9��6Kt��q{�>�=I�����Me�39iQC,�����>�;�Vc;��f�����FI�����VH�5)d����$�N�4�2��фj�!b�Kޝs>�*���g���y�\r��ضF)Ҝp��N%���:�[@�zG�n�,�#2��|�!?\����NGǊ#����(%���Mo��@\�ʱ�iIa)�u|˿�kW�4K��l����1&�(�;`�:�t�V`u��P�f���t�0��sܪ��|�VŁ|-Kq:X�Ƙ�fC�B�Y��� T	�/�[�&�硅~���o�0&�q��f4��8+r�\��ˏ>RI�2��zYjt]����z78h��!��5��p�����8�M�+W:.4���b��_7�z,�g1R�B3�Vm'g��䕰$��[�rJ�5�I�N�SB��v4Ӌ�h�=��{Z�����`珿�]/�t|z�Y��Qِ��a��Ro�������.��?j��ؒm�	����m��ۨZF|�R�Ƭ��H�؏����6,�7�G�J�q�Hn�/�V;�G�i�@o
s t9����'����Q�ݮ��6ND���Fs -�c�Q��-!r��*]�p�NH!k�ġ[��ý5���8��St�;l=V*蟤��X�9_�,�]���L/��d�A���v��ʜj)���9T�L���}��f�&s�Q��H�	�޾���β��U��`̭o)3;Zya�;\sg7{��zm�b�N}�󘅌8��'�6�����88<Gz�R(N� ��>1Z����jjܝ��[�H\T�^'�*>�ֺ�^y��J%3d��!,:<Aף{��e�g�\ldgj�3Z��
����k�	j@�3Ki�Cs(�}i�T����d��{��)��R
��)��n���%p�{>5h|>(_��Cp��0i �D���vS/��/��jf��,�����m��,�Εp�;�RL�ӄu.�eY.�q�ɻ�]��F
�w����m�$n��zP���rM�C� ��GYX_����I;$���H����% ��S⮤����l�ŁSýL���@�57���eP�h3�����V���� �בC����^���Kp./C�>R.�"�$4�>XG;Fy=����a�]^��Q�x�����N�Se[����Bv"SE��%�eL�����|�E�6Q�s��
������?a����e<I��I�<��酌v����̪����ep���yxP����^�����e��H��LB���"rꌳ��ۅl"�*fZ�1GW�ñ�?>S_���.����_Ϗ�Qp0Z����1��-���׊�40K��p���d��#�vu�C"���R�Y��sW����k�(_�?�U���������Jج�^�$8|!>�(`�/	/9U�,�����w��� `���c��@��&�+y���ʏ�\�w=���;U� �Nֺ&�8��z�i���+o�"_p�r喊��q�?@b��g�[F���J/	�c��%�Y#���[����X�w)��O���a�2Ư����Њ�F� �詖���3%���V$g`�����qUo}p�Y"�E�\���Z���m�V���J��츷�}2wI��Gu�5���'�5#b���%T��Y�S��W��莵���S#E)��
���p�O�F)�'������ �ڌ3�u�]�����~��M��vN�Ф,�(��Ï0���;~��d�du��`j�G�$Ywk��
�����3�Ǿ^�6��<����5�َ���$��ADN[(�:����=��4��]�����m�m5Pj�B����tgk*�i%A�DC�y��x��Us;�����B��n0���kN����A�Ŝ4�!%�1eZ����!Z��E���q�>�t����������k�pm@Z�N@����ךc��H#��:3όف�p�-����k���>؃����D�k�1{n>;�/g�,�\cb��5s�G�i�B���_+h��	����ބ�6�����G�b����(�	8 u���lDԦ�4�R�;�#����T�I^��'ݑeWP`�~
K��!YU�jx�e��Ss�8�o���]~=��N�Ū���D�X�Á�L�C����`�n5���~��,�qn��&W^�EJ`�������q���uyf�;�)@�9�TtY���k/�e�K�E�JŶ��āɂ?�]�c�5��3R!�*�Z����v�����Xe9���}����IΈ�Q6oR�lx�|�<���ښ1=� ��L�k"����/ʧ�U�!{Z��=(f1����6����$��0���Mx��s&(��נy7X�Fr�2@���R�����8�w_/v��v��#�0�G�kM�=)oO�$�@�A�>�Z�%����ٹ�^���fJx��9v�Q����ғf瞅-)������^0Y���Yd�6�x�<3vR	�=� �
A�����S��z i�Ӗ�VgXƯ[�֙��&���[�A�$o^n�w��q�n�j��T��;�	Fж��Z���i0$�����JYC+}����掗׹���I���h�������̄�rގݣ��@�Y *�/`=�<��b��nP�g�=�?b̶�b��c=7�9�����Unu�G ��X�X� 0���N�tC(Ӄ�����n&��9��$׳R5�"��y5�{}�;
H�E��q�xA�T�u��ԃ��B�ǐW\�Hĭȱ��7JJ�?���{���O٨e!~&�"���O$�O�L�(��j���Χ!�y/L� ���E�2�Ή�	�D��چ4o��a��U�-�Pf�S�H����q6f��E�U��z sNmmv�*�2$*��� 6���M'���T�b�^3��d��ֶ��(ј���*�D,��>:��fet�$�������&kɇS�[Ck�8�������ǅІ�� y�3�n��36h�����v=?���iA��K��g���ARL78&`��B��܏�.�6}��D���0�r)��@���8�b��v5Ꝅ��v]~�h.م14��j�#�Q��w��w�u>�0�Ŏ>FE��/��Ϥ�W��S�{��1�si�@�u�/]���oƅ����x啐�zy�z��e�4�/r�}|3�.%S������x<H�ލk�zR[:�S���XP����G7"��N�V�
���X�O$��I��Z�ĝyL6L���mh����/ז*Kd���N��'�RDᾔ�9���%�f��t,g�p�W���0V�.�&s����E�7aq�Uʩ���$�M�-���T���N���R�a7{��t��6���!�`����i�oE�x������^l�'p��ߎ[������'b�L^�E�L�&�,=��Q������Z_�w��V�,����E�)5�ۑG�ܼ�+
��&a^2�c���!=*G���~�:�X�H�9d�F���7ս�l+,ެtK,ba�����	��MF�l�
4�-�!��bQ�� *�)a��aJ���2#��s(�(��Sv0��l	ȁ�P�Ц�E�7$k6�{u��Z�)��������zX���O7��&��[���v��B^�JO�P��i��6����=��E*�cG����_;�|��dov�<��k�I��vRq�2�Sn�`�C�2W�o&�N��@q[=���H}��|f�q���|.+Zw�_?�g+���*œ�V�Q�;�3�q��g�v?~�Ze��쫐�A5��dd|�G�E�͘����M���8E`�7~�f44���7�alS��l��x��!Ьɒ���f/�=���CkW�<��-JH�W͚����z� {G�m1����<8���«!E��&6�6���4?,�n@��Ç��b�x�Zf�r�բ���2@�x~s=���i١>�y��T�\ ~��u��F�Ǌ�ؑ��t�Ώ�$��e$�;������#��O[IK��؎��Z�û�c�cD�;�f��h;0���=�I�*����K^W��l�F�������y(�,!���L�`!J��w�D���Ù�M:�~�b����LxA۞u�H�:ikoe;I��pm`h�X��T����q��l��<S�j�|����e��ȥ���	�&~@f�V�jn��Cw˝&C"2�5��Xߵ���
WId��y㿑~�WYu�����r�Y��:ֆ��'O>����}��/ޚEsX/��Q �G��`j�yx�^�Cr��,�+�Nc��Rpa*Sa��G���SI�a7§m��� ���%Z�ZlT��:��7g���6
q�+�lc��]ԘQ�~o��R=��p�z<���U*Act�	玔3ge��j��&�_襦7�i-�0���R��R&�u�����B<�e@΅�!�_Z>��#+��{�h�k��/a�峦9.q3-�Ŋ�������I���|}Xq�ް�	�49II�T�y�3�/U���ī��K���|J�R�#uܻEՆ��8�2����
�?1v��e��7�t����^į6���W��_A��C"��z��o�<�+�9�Z�Z���zѨ��a��k��XҢ��R;��~��?�o�H㏄�'�V������`�� ;P�\sd�R�U�@�9�I�&J�)�~E���ڮC���
i���%g�OP��|6�?,���!ZO��-cϜ��2F����{rmԅH���20l��K�l)4(�Y"�+�G�Yɠ����h�g��y��kV4�'۳�&��f��������j|ɥ�xJaV���1d�׭�������2���7��6�X�Bq�-�0�R�̄�C3x�8�ԯy��E)mŊ�~3h�~L��Lř4�L
�0�n�gM�2�{2��~�9▃��g�����Uf�Kp*d|�/̆Mv��b��}n��M0�$v�lq?H�x�"��&�+�v�?&eߜ�b�`�֚A�+f"%��ϴ(�*}d.%A��w^������L���Np� u�/U�wK��F�^�~	�ǁ�̔�t�z�gy��]I�1M��%џ�/�qs-ܽn��{I�a)�~���:��J�CYh����J�H0� He0��u��D(/�i�c7��"Uw�|Q�e^����(���xu���3�ڿ�k��7��ۗl,=*Q�&�˅���\8]�]M:G<�n��P�`OC��&/��	k{mc����|}V.��_��'�.�(o�BuͶ��J�o�+#=I[S ���2�3��W3�K�RxEI�FL��鄖d�L�PL;����J&��{�+��������FZ�,t����1�HkJ���c�1��_�,��J<����_�)3
h# e|,TE�����5�
����|[���T:����'|7���ķd�p@�d�fr�N�1A?U���0z3���D_�/�4��L0����N�޹��dE�bQ/�Hf�C|~H���*0�Ў��cN65$�<�Mֺs�F��A�?��z(H��pp=�Zo�p~�{���9��45|u(�#ힱ�j�:x�x�Z!#K?0�^QA�� �c
��n��De�J�d	�r�k_&�v�@�)��^��R����Tx�9>�@�۞��g�y$w
Ux�ᖲ��ka�����`օ�N����~�a|V6�����:�nb�|�8���D[�2^�x��=%HD���rZ��bR�w�Bo�q�ՍiL�#+@Yx�z8�@ 9J��}+��[�s��pZ"�)P�b��d�ͩ!���x��{7 �FG�¾J|"tS�ؒ�*8��c�7VR*O�
�
:�vА�C��G��ю0�m;^��2I�,�>B_�7���S�^c�v��=7�,\x� Y�+n�#������������L��$N�$[nҝ��'A�����GQ!u���U�MNe
쒝M8�[�,��N0!Z[��{X��+���\+�'E�=z᫣"��g��%��IXE���P͑��'#G+��9�p�4`�{L8�LQZܳ6���H';:_r�D�Σ�3ۙ�������=�rІ�[�|2�*�V-q��m�h���%5[�������z�"�6y`���#�%�U�m��Z��?d}�j+f�ZY�ԋ
Ĭ����0Z�G�JX��Q�����?4�������ޑ�@��3�Ǫ�<�tU��|�b;��'�O���X0�͙����9n[(R�Ah�!���N�N��o(���?k�2/�b�L��b5*BU�ٓJ+��A�A^#-fY���@&t�
\��I�Z���5�����$&`t�p�����
��&�,Q"�n�l��y�y��i��[h�3�qOI�3�Q\Ŗ��@�aɟ�N�r�>H����G�rO��90$A��*���?,.]��Q�&�ڒ��z��)�\�#ez�ni��� J��61�v�U�
�'Ô\�}�>S�b4����f��2%�xF>�����\�;�]�%qa�T��E������A���~�!D�籅sFt�Ȕi$�����Pvh�Ků�V����a�#O��_�|�$.`Z��qs|��n��M�3g���H��c{�u��S[X$k
����{�g��������m
��a�f��ʀw��stOad&��P�{�G��d�flK\=u��^M�-J@�a��Z���Ͼ�?�q�!⊣%m������P�"ˤ�ʹ�5�hJ��S��u��f�����'r�����*�-5=�ME�����˟���BVU6���o�H�_�?�{ ��l@��	�>��[���x���\ա�/�wN���^���S6\��y2/�vc�1���q��4�xdf4u�<i�o5�5k�#����R��w��.{j�۠>;˔�� �Y���pU�U������a6��M�H=n�lTM��K�〓_My����)Н��Đ6	��������
�qz�OG��"��'!w���&7�m�hm0�S� �u#��K��Q���T]@��̖)�(vn��10{�g��Ӥ�}~�d�='� =�ܮ��Q�޸���U��	��e��ޓ@_� �~̯K�n˃D�a<q��?f��Mx;����R|�,�ʗ��Ok(� j
ď�<t�a�w#�Q��i�0or���"�^u;�	I|Wz�ģ��D���z����C�����V�6�&·�|�/E��t��.���
���n,m���^;B91���"�$4ڦ}��-�4sh��o�e��r���%ѹ��;�58��/2��d�|�jܐ�Q����-Vu��8ȡ�׹��6}UO�8��n�:��괵���y�_�`�#�Z'�8|#�{����?-VF�)���ロ+!N�����j۠����=�~�j��Y��-��I��HxY��腶Yc"�js���7�%_{�y
�0Y���~gJ �l�q�2}�m��� L� ų
�QC�[M��z>;Q�H�X0�AzNj46�X0/<��d�Rq}�D'�vҡ]���(+
Wa$V���"de�)��@\8� �X�]�+�u��ל{UV��}��?�(9lឆ;�qp�f�wS�r;=�=dK�Y��0�c��B��n_�Q�>�3���'�)ł�0���~��l���D:��	�U '*q�����f�������ZU��^u<���A������[R���=˨�aώ���c�3u��\�����>���'q�0��mǘ�e)� ?�w��'$)Xt]ѥp����mS��������!��
l�y䏾ʝ!�ٷ����X�i �o�.�����?ޣB=T 8G�}�Rq>�d\��T�^��;g����Y��{p����ӹ�(�-Hk��)G�?�"�ݡҠ2I���[�����6;G,s�a�.�Ջ`�����Kt魘rl_�����%�Q�z��L�Px��`�����E>���>���}25a�t`�6t3��^'�T�i��2������+�j6;������C��O����j��Zv�;���<�U�ݘ�p���bP�_�ʂ�#�:�>��kR���[�2��Z!ƀ(zz,Ow4"O��hᖆ�>>"��p(�f6����
T�^�t�4�\[�S8�{��rQ��p&�A<}�o,Z�D_sÁt��ccapZ/)�,Y��gٯÈ>P����p��@o�ܒ+��?d�F�̻��&��<X�LL0Y�&�d�UČy�S�̀��۱N%�,>���r�/ʪc�E�O=�'d0���9���7���g�D�_��;�Q�2��f�T@��qcM��=[a�m��B{�nV�Ӥ���K
�Y������� `��y�����]�g���B	��&�	�G?ȵ�i�t��p3!	V�,uc��\㐑��Mutأ8gϚ�m����N���mz$��i��ǌL��y�4�w��w���_[���oa:D����w0��9Ȕ��w�[ON���I�i���>�O())�-8�k�XӀ7�,�W��mQk�f�^����d-F�?���r1h��y`��q�v��-U�*T��ۓ�d�����U`l�@.z���.�lE�Y��������}d�v�4�]�C�.��(J�"��v��?��}.�Ħ�g�{Z����[�^�0�R�.�܈�}^�3���{�$H�7���-j2~��U��֯�c7v�Zq]��ш�Jjk}����qē�aʯ�`^�i�ҹ���x�ݪ��� �͙[+�"$๪V��}�,z��<�kO�׊n���?����._�'����h��.4�`K{�T>�����_����j"1������H�"g����[�%	�-�xo����~]X�CEz�zP���&��#��C�kK��� ��Cs�_��j"���#��U1(�7�f�d��ӥ�`ɯ�3 a��s~�K��֛�+�}3���E�8�V�M"�UB���A�.n�,J��h�<�>��d�9|/f|��G�%��⺌!��������N�������p��c}u���s��� '\9|�m�[k�iԞ;��"�
��1-�v�tNKwRI�5c]�����b�u�E��������A���G��V�^�t��^�%�	[O�9����Ƅ}�м��J��P��L]DJ"���Ƃ�j^LX�F���?���P�R�5X�PB��1;�h2B�������Ą=0è\�j.����0,��%Y��潥��e2ٷ4(3�ȕ
�l����:~���;L(��	��q�nP��Ѽ���-��t��a��z#�LDJƻ����*�Ʉ՚i=t�؛����xT�u(os8EP?�T$Υ�$W�������T�.�"��!�*ތ>�Va.Z}8R��YK���1�Z�,?>�m���ϣg��{^ ��ù��.�#�Pb���ˍײ`��G��9̹�����^����bfC&�Z�-_eP��ܲ{��D��y��22�X$��Z������u2Ӛ�g���n�9	�fx#�}��1&U��7��|_��FB � c��a#oE9\�0�jB?3���*6��;�f:�Pf���2��?WgH���� mE�#��.���YΊ6�E��w�e���M-{��N&�����c�)gsM<4~�><?w-��mK��6,��T~A�^p�V�ϤC9"�Q��>c��"�5�8�L����B�
A�/�f����n,'�+o�Яp��n#j ��h�Cp�D+D��bQ�ޠ��HPs�ʖ��"c"���qc+�j���p�u��1.�;d��P���廫���L7�4��Cas�q�=��&�|��pV��癕-��O�|��߲����A�'g��Y?i�����p�i*�c/ܠ���^��	7H�m�k8���c����?Cmu|E�{,&y���I�Q�eV�9�D�o�G�t0�p��,������TJ&{��W��@ږ%��W����n��?'��B���	s��dH��-����.�P5wߊ��	��d5σ� �d�%���=�u(��k>��%�a׸j	�^B��r!���*��/�	:,J�������-(�]e�*5�z���r�v �'�,��ɂc^�:��x��+�$�mݴS�Ǜ$;�����	�n������1i`;q�S���	�ƶM=�5Ͱ�|t��X�������4Wl��:�u:#���Н?�!;	e��cHc��Z�����"���Dv�2��8]�0f�@;��V�N�=./�M��L�D�'�y(d_^'w�b�ؼ�y1��U�
Lkp
E�Z�l��$�軥���|�V��Z��{��!�1�̥��#���w>���_�W6e�61'��$����}<��&�/&��و	jB�q"�'v��i+=wL��[�y�Y��7q�}5e�Jh�w�I��=�hBZ�>Gj����G��l�aG��D����!��z��%lGm����>�T�����L�q�=l���Z�Պ@u��Ȇd���8�_G0>��qƕ��@~���_؁���\SVC�Hi�h��p���K=M3R��\��q�Y+��+zf<��FܿJV�[�Txx��������u�6�B����Q2���i}Xi����i�jy+�A�^�ePbA��S�l[%9�nTPrR�9�����/Ȣ1 �Oh��rF)ג��P;t�A�tc�\��Տ��2��
QШ��e�&�4���Ud�C����9�g�`{b�����>�1�򤁅�L�k���!���O*��0�;z�=�b1�J�<�i-)̈́Z�&���̇�0h�7�fV�N^m}�J3�L�������βǢƂqN��Qn���Ս	�D�Jߍmڹ�1�e�Ɇ�d��"*�)Z:���v���t�mŘ`|��O� ��=�'B_�8�}�6�Fh�b�G1j"��J��t�-!I3���NPsR�{cg᝶3U2�w��e����\L�8�r�����f��h��*Q��\�H���3(�O�7]s�� ����I��RX�:����nS|�?�1u�I�a�����)��Z��\a�������r��f��B�n�Οr`73�~Ĝ)�Q(�1y3���@o�'�f����z�H@T�H����E����*z�D��i���q�3�𸯒�
�OU�WYJ˝��:�8b��C ��pgkx��x뱍3������~������4��.�MOɈz�ΎEH,vw���ܭO��z�l�]�5�W�ւ�X�����1mϚ�Ų0�R����S+z����>��@S�v'\k4<��HC�|>�����P�[[����7�p�u?d�$��y�R���ת��nJs� ��AJ�Ǣ@抑�˸8�S��5Ȥ��	�ik�G��7*���C%hY�;0p�w�����у�g��I$ ����_b
�����Hc�?q��˗����&�IժD���MJ?=�AS���q��+G!69玒	�\�	���z�M}��G����q[uL���\���7��f��v���\zݦ����N������K�Ϛ�H�����v���I �d�'"w���Π�kc(w��'f�Ga���I,![.�q�tX^R��"~î��P�nHZW��p<��Ab&{�7�+ gdgy�_%|Й�nF;#5��&L
5�Qb�VQ������CԚ6�O�~�`���^�n)�F�P}7;*�L%];�Q�	�=��ϒ�� W�3Z����)_@.� ?&�� ����"�.����e�]�/�3�@��<R#�lx���$��S`|��o"�)�K�}�y�J�>�'>]�Il�&��)R�:�t;���+i��cC�FQ��{��ldw��m�vZɐ�����Q�����*+!6�z5���5�7����C�������b�30�N��3�.D�|�w	j��M�	�gLl��k]đe�Y0\*Ө@�.�åzi����`��pN��]m\�c�f%w�ױ�;��&��σ��?�"6��2b�#\�:��l�G�"��s($Nx��)�9��iE8-V(.ii��~�N��B�P�Y�T�`�K]���׋�Z�2՜�9��-�J��b騴q�@^6�Ǭ=%
)��	�*��R�[C��4�)5F�Qv4P����R�r������[c�Ĥ!��Nt�q�(K��tnpY�m����H:�,8�����Ӳf"�vj�d��_
�����h��D�1͚�����3�b����%��X���� s�����e���-�|<�X�>�J��Ht�a*Oq������b2�<v�	�O'"���ӱ��0�;��y>oF�nby��	���L��ͷ>ײ�XJ�<�{,Ue�iK��L�H���D�2�
E���x[3�+�H���Y�	���(�3[�u�@���`B�2��B���H S���ſ2���I�m�|M_�нB��J���4��O��ȥ�tG�G��#�VR�q���v��~R]�+"7r�ѧ�$�1"q�t���_'ߢ6�Zr�h�~�[
�Ĺ��|��J7�,�px�c�7OW4��`��^sf�nة�,���g|�z�\�4#VPa:qҐ���wV��,��y�F����2�6��J��Mp�]'�9�x.r�f��U��\u�z�a�d1�3TM
b2dƍ ��_X%��UT2����*�@6Az%�9G;X��<8ti�9��$�l�+H��|G ��`0|��
V���:��^��4P����� �y�����c�s������H���!B}��l�n�c�]2���o@��Pv�G���	!�.p�0�r�dՋ�&ǌR~U6�9C��0�Z��k�]ʇà���������SB�Ku���43�ɵR9b*����i*�݁��+��@S`�#.��:�(0����d�Go}�ݒ��FUP+��z�O���U�=��7K
���y��ϔ=��} ����=�[��n�u��6��g�ü���Uf8 ��"��"�����}1��`p@��,�.���&I��_�c�eQ-0P8X��}�_�<�2�{��T�;��1�N����o����YYr�y�6>��R�N.�����Vç��jk�����=s\o8'�a��-'����R���{
!�S���W���k����i2�bZ�����������$���� ~�O��M9?��V���G��b�	�ԙ�{)�Z;� ��h�X�4%�De���$�$��(�6MBX�!��uJC��/@*V(yB"QJ8�����e>,Ef �HZ>�K�u��6�[W�=|c_�*�kx��}��s�fn�~�&��t"�	d�A��։�NC��:��I���0��k�����^��7��>~��1m�eS�����jm�Ǎ�{X��y_'����W�J��UR���k�}(ǡ�2�έn���F ��_ᏁG����{��]��@K���t��r��d��\�]���taǹR�P�{9�`y��|���٢	����;Mim����M���P#+-�0�Y'�i����$�<����@RXj�D�"�{��]�oR���3S��2�cʻ���Y�7�_k�4i6_җM7��*�=rm�V������\?�=S�j5N�o�ڰ�;#?�~��	>�%�z��m�K�<���aZs�\toK�G�5�{/�E�B!)���=��2P6�,Ma�+�{m4���A�{��K�W��ۤ���.ߚ�%-��|B�#�n��2�F�O�H\�"�Yl��6��.*�y�M��Y0��I�c$A�nF&�O{唹�8u���Z}۩�vz��z�p~E��Z���q�C�M|U�:O�*��͔�o$�k
�L��=�	6~8n��_nC��6��.�ψ�+�^l|�\L�G3H�;�Pa&�Y�ض&!�d�M�c�~�!���艁��[�����E�H�繳#��$��p|+x��k�����y^�3
���{���X���q]G����ӎw=1	���8u_��J~��R#a���c_���9 ��s��+��a:������mڋ�ȡ�f&�,�G���}�%���u��Jx*:#*�g]���B���	�?�3Jm,�Z�@�>�C�+�5����5� @�vR�[�<�-;O4.yЗh1�:��1U��F�-^c �2�S�<�km$aaN.����@���
���׉��A�!Fp?�
�Cp$���,�!�C)�ƌJYVN�KHX�4��[/��$ڲ�;h�Y��(.���/PչY���)�+���2����`���������\��u�t�|W�V��W!D`��-;s������q��F��@�[�`�#7y�$C�ӡ/.��(s�m��0���`MBXǗd^O��?4L��/�0����>��R�CdT�w��P􂗤ʽ�#����h�a��r���_đBI�2�4�+GȌ��a�$�D2���&=6!J]��z��z1�J�%�)��������EDY�c�hI���J ޻��د�G�jч����@�J7�
�Hf��JPE(�-e7I:�U��6���K��j�Y��{�ȯ��-˻C[�#��Ø�N�c�~�9s�]�za2z��E����c�F�H[{��8�w[&3+��x�;�>ɣ}!����U� !hg�2�z�ң|���̼��Ԛ���s����d)�����;���~�
�Q��'�y����`����C]�(�ڪ�L��� �E�� lW����W�"7� ��XCn����iL��+�F��ɼ8T�G 	\2� ȋub�w�*�ɍZB��rW���<�Bq���@4��~���We�5!A��CT��]~)�D^�SI.�� JC�d����4�&=ƞvb�Vq���� ���ԋ��v��0؁�䋢��ށ��t?/�~	v��r���	Fl����b�{E^�(N�%�Τ=�$m��{㺌�m�&�lJ���	۸ԟW�鲽֛w�n��Q^�!�H�MO�,�_��u�i���(ϝ?�>|�}��^��ޱ"O�.Z��?Ʌ��6ml��<O"7���렁�E\_GTS��������^�ۧ���|�D��krw�<m�Ѕ$N��,a�ςw��#�l�s�E��O�y�S8�����PW���c��
�H�p�XX
�G��p�;�Pa��b����!��A�᪅H"�d�3-�+V��w۾ًic��u�=h�֙�����0#56��1�A����� �/�.j�3���O =��d5|�L�
C��"i�g���c�!*�Ƿ�7�n���N*.������r����_�Fk��&d��É
�'*v��Z��d{b7�;�(� �Ԓ�vL�jS<��o�MM:����X*q)�%���[��@���N(�Ȏ\��}�<�5��p��W��e1c��	p!���Ф����d�키AB���|�ׄR�;g�%�U!L�~.���Ĺ�)/�-��X#��g�k&�^Ȧ���Iy5��'���,�PLIh>��hfJ�:�}߲C���_&>�e�+| �����>皔�:7-5:r@�<AnL��S�ѓ�Jw�u��f4�t��8�8�3�PQ�����FP�G�zM|:'�{���KJ����b^"���N�7���zǬȭRO����p�R]<�(5�W�<�����o,������q`1p�y�Az/aCq�����@�\�@
f^5]�8W�a�����f�� �o���	p�K�2HM8��:KՄ��t�!%�a������l�,�������ݼS/�%r�QXj���II��&/��Ŷ|:�o�S��^�_d���d����M�-UJ���g=#��{�i�$�ڟ<_]�ll�f�v�pH���,S1��'���B��5,�`�S$�������@nm7��@F\��9�=R�9SR���XWEK��UV�(J}�:~��X��1m�4@tyV��I&B���T��+83J8@9�S��	!���A޽�ǕF��h�@�|'f�|�NnL��Kd��A,v���!�[��UbɧT�2H��U\��9P�$��(d�ح�X��^,�Mf���fG`�;�A����c\��US*)n��(>�0�"
^Y �/U�y�uh��L0�O��ީ��"����kU.ÞPA�%�*�|���g'n.�G,Sx������tJj��,�\����G�������%�������ء)�9�ύQ�b�zu;���pb{)�^h)�*-8΀�J��09��¿�@��y��'A�P�mR�_�5��I�ֈI阑�`U��A�>q��(�� �;V0ȟ�Ci���Q8�xJ�=h
������bN�� ���n�H��5j���]%N��U8�!�K=��a����Zu��Ʈ�	cTB��P���5�w����/'��j|�e��[��/���d�9d�R�2*�`3`�̐N|ן|��zM�����������G#�c]l�bʶ�(�\��ﬃP�ۂ*����@J�!�5�9d��SvJY�脄�,��T^J�����a��[�f�)84q���kt��K�$"<v�f� �C��=��SG�a�P��!DgD��c'3�Ek��a�u5*���S��'[��11aUuV��׃��-�I��"��1���/m�S���$l+��@,>�;e��/U��j�h�8 �����D��꧵��r#�?*[��7���*��L�S�|�^�?�q+�p�p>MַhI�r��>�i�&�I���"�>Cׁ}�h��a�K��B��_�Ɖo����k�nn?
�PEQ�*��EY�v�����S��R �e;p��ů�[Q�ڜ�-C�7��JW��æ��48;^�{!+����%N���W|o�#eΜ�ݢ�5�"�U�)�)�W���B�4�"ћ���=x���=E�%��~�A�����j��z��2�P����Y�Į_UOռʿp�i�۫ɀDSj��o������ZF�A�E��RW~�}O�	ش(����'j���u�3�i��߈���U�q��t��@5�sk�M�F�pc}0:�u�|a�bQ�mnQ�I-}dn[#�x*o�G ��M%�FeN�Oi��L8��ф<�z�0hC���:\�bC<qd���P�(|
��3#�n�(I�Dw��g=_+����& 	NC{K<G��J�h�+%J�vE�H�zhg��qp�����W�86�����雼)Gƣ1�K�ށ���J���qI����XW<�NV��'&"w*T��� �����v�V���R���6����Ω�:FM�~ٜ\]�l+�`d�
ce5#p }OV�D��U�ZCLA�}��qh��:����������[e��vb(k�t�/*�{�a�%��Z��s-b�����l����(�v����D��F�z�+�.cѡFD��
0���@����u^X;�L堻,=}�d��;c�j�km�g:�K2�v��c�(mξe[8��(�K�N>RV�����j#K^#�ȁ��aDP�d�����v�����D�
��>�e�����oV�Su[Yfx�ܿ�\�K����(��l���B�5�E}r�Y�al&PvX�b��O.���m���X�����^�ǉ!!Ҕ�R�� �JP��V�<Dە�D�7�c ~��$s�c���*<��T}��UP\@���Ҁ��c��/�E�|�����������s�.�F��F�t<�Q��%���Ӓ�R�G��d����B&-�!�->[�:%g���l��آ�(����_4�ِ�>�r`C�7N.G�to�V���X�9�oo�^Lxc���؇��חqP7��2ͨ4ۦƺ]�g�A��u��mMv���{.�� �L�t�9l�T:�ӃӞ`��'x���쏉N���Q��������6��S�.J�	y W��<I�E��][G-X�6��2�7�~[/��f���A��,�<&�/`��=VdZ�C�����(���VȂ1�W�x¹ly�o	{l���8&�*�&��\�F�`2=0&��G��i�$@�Jʄ줕��5��B+ �A~����cG�P�FB��f"w'���pN]1��~<1d��(����z��F�Wc��"ec���SEJ��e|��|�aZ׉�mXI��*z̍y��B\��>�"&6�	J�wZ.���l)>($�=�E��$c�h���f-�R��� �=��kq���n��f����qĞ�l�j�����fdeJ�:X�,��|U8m�پ|�a�cG�?�=���Y��ч��KsT�o�C-SX�8��ѯ8�����)g�Ԣ��	�z���&[J�R��6�������?!|r��/�UڨW�C)_���\��G����_�H�UL��2_���`X<(l��R�z��Y�9� �\ԝ[�i�)t��\6"��Q�v��w�FcϺ��~S�L�ɠa<aS{&t�E��gȳ�GK�T���<�����:�LvG�DfV	
[�g�������9��D^���CX�o��A��4�&�Ŋ�q�IB3$�D>�3�N1���_����a:�]h2�d}]&��:�F����E1�K�l:]:�K"��b�5�.�ܵU�v���ЀR���w�aA��c�ۖ��J��h�M�Hm'w�~���Wp�U�-������ҧ�qO��أ�E�S�Oo��xT�!�K��H��17�-?#�z�r��m�w0���BJ�Z4lh��~W�RP���H�/R?�輥܅2��x�݊{;����[D�;L&Tǐ��(*n���|e�
Ӏvǘ��Sܧ{Kv)��~�ul���t3��>���ԛ����W����;���=�;j{E���P87���IX�^�Q�*��bH�s�&���¥�1���TK{2�MTz�q�h��X�D�uR��hhP��`�ct�͋�$5��Q+'�7�|G+��,$P���\��y�&ŚZܳ�ws?Yư&)Z�BC�gv��� �p*�3~�\Y���{#͋W��FW-�����io�\)��/xؔ�����MtkI�y�$�CO7�X�H��u�����ґ�N�I�]����n����kT�,�
G�O!��/g�����)�ө�Q�Ӻl��	N m� "i�Z�"�ض͙��R]����u���-"x�hvx��h<���i�O{�>��V��i��f��F	%9M��v�| ��B�.����S�e;������xn�6�s�=���WL{�7��@s��ϵ�1�{,�`�I��'
�#�h���F��>��6�p6�4p �"7�h�azn���?�`�Iao�|�k���4��֚_�M�;tR���T��+��I�\���e�
aB�~×$%jϏ�������t3]�W͕���}� �U��X�&��[�ē��7^UeQ���;��t�4�l�&�>J�<2s�Kt��O��3&���#=P��=�`:�F2�p&�׊5R�_��Н��K�bN���,���kK��`t��xa�«�f�g���g�>~�kȿ�j�C*��Ǳ��Q)� �x)cs?��,vݲ�YB�)���H{����m�=�jMM��s~,�"A��9�?���C���?��������P0���Хi����
�+h��G�LP鯒ZoS�&�؟�OR��`�u^b�s
%-��<��0��Q��nn��d�T��p�O��+���{<n����zo�}l6��A���ذ�ϊ��{Kl�7F�S��T	0�@�%'|\z\ẑ�a�I��ă�Bϳ�ɬ5
�k�f�ET�}#h]��S�������g�|Ype��Yo-`���?���=����d�ߦ
L�����KN�4g�i�ʣw֖97������0�vXL���L��[v�9�S�@|�I��Uk��4��h�}ғ���@H�>\� A��~���sNN,X��]� ��]�R��	���5�Vw�_����	���Н4guS��2i=�9�0�{�.ޛy�g���I$)�*�H�w#�)��k� ���C�Y:I�h�ߔ�=&���U����J�aӎo5s�Y����p8�*Oi!���j�~)�S%�n;��M�
i��"�a���־*�	���q�c(_��u������a1`�#]/{�D'�Uf�_8�mN��2����U������M����ǖ��
;h a��Cٛ�;WK���U�1��F�j���D�vv�Ŋ���$��j��k)?��4#>AE���ե��]�'�p�˖jCn1��o������VZfb@�%��1��ꂐ�Y��i�2���n��<S��H�\(W��\�1�^��/��ʏ^U�y4M�F>�80RR�A+0hԛ�)i���~#22$X.=.�����-X�^a�.]��l�8�;��0v`�07�I7�ӱN�����N�F�pl���ş�fVt�e��:�:�1�<�iB��]Jq��l ��|���C��lHW6��5�5�!д���^T}�������j���&<Xc����3�����,��&u;TY�𴪨�f.qf*�pv��$ax�Y��;�;�q��*���q=�����0Dw\@m.�k�	�a����X7���U�ǯ��o�ʒt/�w�;��60#ҫS�ܶ���v���1LbΚ�H{��B��Ɇ4�1�j�
l$'����v����Ւ�mI��.ʹ�.��?n���[G3}�e��n'Je��*�q�_FN�Je;�\k&���[�뫌���i���K�K�wYp���"�-� � ����J��,�J�2����EW���F,i��q�sQ�e��ipq$��c,�4�M��|c��%I�C�t��`wI�+�ϔ�%�,�6�}��L�k�� ����+Lh�5sʕ�G��#m��t��cx�"?i"��y'Of�;^��P�m����a���'$hD��h���A�z���m�l�F�6�Z.&��3�
׫��Ɇx������E3/Z����v
�t(I���}4�:G�I�>0[ A�̱Z�@/����~������'���LI�_b3Y��	�/Ƣg5Wɰ�8N��� ��G?������<�Ut]�= )8���;7���Sf��1�\p?��K��3"�����Dh���Dr�x>v@��̹�C�ĲRZ��hj�"����AX�����!�008���/Lk�B�-�Ag�dpRu��g��䗮L#=��w��6]�3����O���2�KtTʶ<W�R�'K��:���Eh�� H�}����Y㮞t٦+�&Y���_A�;�#�z�49�jײ��o*��J	�� '��3�d���.D	��VϹ�i|5���}���YEэ�~�ݏ��RU-%�ȅ��T�L����k�.�4��>� lǻ-$Η����3��~J�'��2PP��.M��H�2HƉ�,KX�)��S\�F�'68.Z���Ms}� ����gbcfR�($]T�Ƌi��U��e�C���Цǡ��I��mܔ1tw��<��^0O�$�(3a�u�Za�h�����4�v�6J$�f;��!+\�� -	o$N���j���â�wo*���n4K+�gaqU�g��rhmv4d
Y�#�)e�h*o���1"�����^Jt�X�����ƈX�}t���/-o�3�2���?��@�9~	ڟP��c��� q��\�z�g�Ҫ�?+\	@@��`'�i5��V-����Hc�v�����*Ԕ2_���W5�T��V�<���fAA��zL�u����O(�c���<j�1u�ܰ�@[f�|�:X�!W;L�*1K-�vT��ּyp7"v���9@FXg�|�+��Uc&P%OZ�v��:�?/�<��"�'=N>���v�d�}/�k����u�i�ls�Ş9�ٲT󩘼i@�}Fس \K���ۋ;݇��E�T�@���zjs���e����F:���=yE.2�ӾF!���n
Ugp��8���5�7f��8;[���a�g��du�٫�\o������A�� 5��멬�?/L�b��^�@��ϐX:��W��"�6c��>c��+)_�.^��`�z�m�ƣ~?��[Be`��HҺ�� �	��e���,�H,uX�VW6�v4��J��u �~�
>d�1��O?�.{�S(|i�d4�TƺI�˵7S,W!��E��"�M|������.'<��b��d<��p�f���3�M���o1�5�����b\��-��z��o�Ǒ���̈́�@����M��{lZ>���sB\������r����H�z�8�5��n� 8|E�+a_�x��	�f�n̮u�_)`��W�݀5� �a�ǩ�@-j�����C(e����8���:ѥ�-0�A����>E��l
�Pj�����~��Z�S�X(���iwW}x�\�����M��� Y��Qw� .�_ �;Z��P���� g�VK�b����
)F4�4��E�D	�vZ-#���kFM���s�r�we�ٸ4(�ꥅh�7X�=�χ�|~��.�M ���b��(�׵�M��.���x�k�h�,~Ye��l���bȩv��I�5�V��q���=�У��qzؑ�Ԧ����1�F*����Mސ���66�G�.dXÑ����S�Z3-/��R\�:��@��^i��p��G�t���W[f4�p�A�r��)������y�E�\	��|��M��ى���ņ��U(�t�U9T��޸f� ��]:�<������#+<�!�Qw���4Y:��"*R{Y���1G�b=_������8d�f�����/g��
���E�{�&��M�^ɗB�~��j��\�8I��H�W� }f����p����]����%�[�a��2��5纈/�Q�-��G��t����&������Ĥ3�Y��lx?8��6K�W#$���q~fj�I��f��@ۥ�C�.h fR��}ۃ�]״mE,=�b6���f�-��O1b�T\_�9 'i�����_Ϲp�C�j��qm�&P /�j��w
7�K�df�i�g`�R'ڽM�'`�%H�����/v������R�/0���<*�P���Z�OWh7�hB8=��<eZ��v)�QJ �ˍ��� %yR_�b]q֤^	g��*Y��<m������2>�y��\�N��@�_�D��])���n�\���U�.��qZ���r���bf�D�|�}�B���(�U��;�fn-+�+����F�A
�.�Q�u�f��^�+ǎ�rI���x/{�2�9����!2`nB+���Ϛ��8!j�>:��Up2l%�3���0�\j���O�%	��~f�@����ǚ�5�XOHRA�c�;7K��fI��z�����^��)H��1��^��Q��*�`�ҟȖx�C�D
��QY8P����JB���.^#=㰨���[�t+����;,LA���������ڤ�{�Uw�Yo�v�oY XC"\�+��X����^�e�g��Aٸb���G�R�ͱ��_Y<�7�3����c&�?a�*�6���y�W�Հ:\���	�t%,2i��?o1��\�ݨ��JRt,?�K��R+az�3��&ŵ���ж-��c6l�;���G@�_�
�5�:�����"�L_�/kwPu�Ow�v'֤�+;��Z��"��C�N�b�E��[K���{�ː!�>+`21��d |䶇� ������8S2�$�.u��']�n�1ة�+ō c�ݴI�����_���S8����u�D���`7��ì�Oph��N�p���(s�a�.~p0����Og��+h�a�����u;�<���Z�o�������)�vA<�҄Ff�+Z���=�Z8�������a�o���{�I\<��\qVw��=� ��Eo��@���\]<7�8���p���3���TW�y��8�����p����?o"��f�o�a̱nT�·��tx��ˌD��>T�.*�rz,Rsç&&S_���%��<FW��o��'ʥ���X薨˩U�YFѾ¡�������4ȳ���/���yWvź��+H�f�R�$U�g{D(pS�3N̥��$���-���M��p��2�)��nP.L��λ�y�˭��������M'�24D;Պw�mvhj���d�I���1���e�L%ӥ�7�_,��m�[����
�,++:��7oM[�ڟ�2Bt?&x�3D,�c�:�vϰ�W�X�|�10
���9��C��hr�~= ^΅U�}�����!S��<��p��%E<�CU�$	��7�ۂ�8*�4�o$�P���h�aAO�L4hA�;��q D7a��K��<4�=*��*�I�C��r��!J��2�A�ۋ��^E�۴�����oή��T���^���;8�Sp� �nx/i\8֊WE��`��Y���u�߉3�M����up�N�����5�
���#}&�K?����	�&����H8l� e�uH5��oj<v����=�*]�"ΎU�cַ�ZhzP�s,r &�����Z�Q�]ʎ+ަf��_l�>&'$S�^��Z�rf�-��~�>�2٭�߼����=�GR6)e�'�nٶ�iڶ��E�1��C��S���H�q �@�RC��X'n+��J��;��\F�&.�{�U��g��~��a���.f�`8̐�S�׶�D����hb �v��f� �����ss�SEw��V��Em�j]�i�F��O����r!HD�I�b�bX�#�+u;$p�7�0�X ��_KQ���LO�C|E�o�&2��: w�}l�����!��ؗ��P	;�1�٤+&�9�CK���k�F����A��ӭ���\��W`���9��S��:PVcAz,l�I~��R�&}[��>��},)��;5�V+���s��]�|63�)�_
����ug��nB��6���CG�_��K�ho	!;�e�5L���!%�Ş��ɴ���{-� �;�B4ޑ-������u�g���Ǡ��>���h���_�H-P<c4���A�k�������"v��n��ܗ]W=F܀���<cqj�'
+/�����10�_��>mx#j�u�\\�H.6��_2!�~�	�����N�j�S�u�29��B�ŕ���L�s��&�kF�@B��GY\n��Q���H��r�(FF 	�����U6L�@Iw�8ᑖ!�h��`V���m)��z�C�ڲ
��UZ{��`p�^K��qdC/r,��,`
���|��l'� ��-n�vv<�=��Я�y��O����q�9*u_��.��ˊ��&��%lHl�VSz�V�!4U��+H��\���1G�1�kpl��IG�������1�\��M��u��2�,Wh�H��~\@�x߇���n3d���7�Z�/�>sh�����>��B�
'�:�ku2������}���?�����FJ`2ɻ�ӿ�a2��ƀc�X�񾬀���TA�v�svxlT&Sm�"�x�L�dg��i�7~���12H;��P<�[��u���o6GΙdu�Q�AO�̓��˳]�,�(ξZ�)�-Yf�-?��y y��\ �b+��#�i»@D����>�ᕘ��2����"� �C��7�b�E��k��O�o������<J\���ߨKf��md���2H8u�<��G�%����?C�k���oyD���!t�އ�����юnZ��ƭ-���BK~�p��?�B��m(�)��>	<h�3E���9����d��mv+|��z��aZ��f?���<��TL�3���x�s	�Ս�VX,�9kr�~��;#x�E�����7j����|���� �%p�ƚ�V֮%j	��@�
b����6���m�8$�s�q�Rr*9v����u2� %�R���z���)�I{�60Cc&6@#'�������1~X!3'�H����%b-�^��3�7��?��q-R�@U�����g3g,0@�w�zH�F���F�lI�#��r��%�~i'�{�M����WMs�t��j�l�IQOZ֗��W�e��B��W@ݼg��~�,ѾC����q��j�"��q�.�p��C 0B�{ ��G��?R"�f�O!%�Vt�5\˷������m`S�VBOj8X��I��K�㏝$Ͷ/C�~�&ADL���/	?�a:���v!�_S8d�����dߣ��Pv��e%EvxN�wÉ/����i����)ZJao�7��̊����Z���d ����?�a�:�����X{sGm�|�&5ɔd�����v�~�'�b-�������8�z�b��?H*a���B��I$���fc�D��7���%K���L+)ǫ��� ��R��(���F�szk(�e��`M��^	�(�p�6����QZ������A�)r�Hn�qxM�Q*�{�Y�S�'�PS�,�0�4�,�|�
���]V�����ۏz�X��)žV�*h掶5�#��UT��<���(TD��]w�)7���'�U��t���<t��F�D¿35Ӭ������z�k�oL3�<Bs�-xL0�Z	V�f���8c�:`���cC����d�Q�"s��X�f*;�g�t�GP������+���y���p*���ڙ�i-IYKZ�e�]�g����.MG:}3��@C�f�-k�1��8zL�t���A���,��C�mi�Q�M���{���q/ӦM3&�&����L
@)Z"�'1tO�R5};����,o�˗-� ���(�E�Ə.�G� 条6h��Y���ģ#����qz�Vsu�l?Z~�Qϲ6J���+�_�d���5w/�26���c������I�������m|���2��'��R^Edb~���r����e��~���7�n��� ��H��-��E5{*�%�h@�(�̈́���D�Hq�|��T��dK̓$D��#�[�NqA��%Y�1�G_��7k:�G b^U���w���%J���-Vk<|���q��iNݚ�$�������ૃ���|��Z���b�%yռH�A�������!C%Z;���C�����o� s�t�u���%l�M�����-|O�d�ڦrN�����Wj��C��o�^]���BLӏ�]ѲF���Q��9j��H��Elf�� H/u*MY}�;*Ƞ�rq��zrI�ȗg{��Yޕ��N�P�{0�eSV�Kp�dnW���r,���V P�Y'����v��
wҩ>H|&���v�Xd6':��u:�ip��h,�!�K�WK�}�AP�cu�����t3aoL��!�>����x/��\�k�:|1�YE /*�>g���`����W���̔+��Z8!���J��+Ձg����^�0dC��.,|�I!૔0��hN�jn��;|���ے�K�
�"�:8U���D ��G������.m �v��;�b�9����� +�)��1�/����k�c+=m���դYZ�?�S���q,�:?������GuǑ7O�ƽ���d�C���v�lO���kƺ�I�vܔ%W� י�迠J�E��Fs��̓�O����0����̰sM���2:q6��j�W�r%���r(�h�fVŭI�j�q�zq��VB��?M���'�%�E"�"qA"��_�+�r��f�?�]����|V��DD�Z�'�g�2�Z�)��{����^��%]�ui�o�YUv"�`eC���Q���$J�/fy��/�-���?Pt�b�B�9�F�o��"��o�O eD5��{��z���B�v�(.�IO���ݳ�;U�ש*���t���y.�G�h/�r���+H�k�B����'';'��2��A�o�TG"����]R�׌Nn��Gr�5����8�6^��;��/0-�����FU��fJ���bk��6"Rp�¨QuP��V`V5�|�Ui���_�G���r}�٣��9�.�j��o
���H�����!���O����z�5�0�����F|��d/37ϔ$�"!�	�v4�؊-���ZF�_���`O�5��B?%��R�:}�@���dp�(�{�E9D1�L�
�Q��)^/�;�(Ñ�Fd����Gt��u��Xb�'!.6����u�(:��W��]*�ݴö�J�$��f//�Ȋ���P�h�uc�o����!���n�������E�9��d�YTy�m�������A�D����)NY�j}�tҿ}�$�f��R,	��e	��hX)3����rGV1��-�`#����6�VK��oz�#���h��l�R�5�I�<2%}��gK�Cz!��.�}0O���KW��������ɁG=��5s�{.d5|N!�I����e����s"���4i昐ۣ\+V8 U������AM�{����
x��F�A��Lx���/#�l�]�)xm v�v�u�E�Fx�MhI���e����i!���$$��� R�QߧΔ��Y_}N�A�M	L+0ޘ���'QƈX/��y��s�@��0�e��
G�%H��L{�|�j��!��%��l/�Q� ��Q���	b��?�}ڴ�G��F�d�Su��tT���@�@X*7���P��FQ\��e�\}�W�Q\�0M�&�އ�)!��|�Qu�x���,�U�c^�M�f�yfi9-d��}��e�;L(M۳���-�b�/�H��3���د���=���jR\T�Li�a�Rc�
��������\����^���kR�e:�e9�L�vvhɏ��]^L���{�'#9�ԏ�����Fl��O)6��"��Y��@�^	wK���Ș�/�|��D���i/}tʍ��M��Qc��/��:�!�^6n-m�}c�
�_�
k3!���c"Z����+�X҄��z0��1|� 7L��1�*�Áv�' ��m�	`T�A@����-p�C6�Kʛ���b�bX��ig�?�T&�'�Tٮ�Q��Ӆ��C6Y=nEd*�g�����4���;[�5ugD�қ9D�Mh���k6su�1y��>�\�	Bm�V.X���������G��v�4o<7��PI/��KY� y�Ln���R@��j�?�e�� I,7p�<j2���mB��x��jA�V	�8�J��(���-���P>��_�Y �q��{J�\�k�~I��9����Ied�x������D�n+�2�F�YRr����_ �����ma4��_N��t����_�χ_�H[劓�3�
\V)>U1	u`����z����3`w��wN��
?�̝u#F�a�����ܑH~)\_�+|�G~��[��GK
Ʉ%�1V�� "N�5̙@����+,��>{�Tc#��Y{�B���,M�g�p�z�1<1 k]��/5�F�#Q����,�>�?�����Л�~!��$�<�P��r"0+�N�c�az��x�>z�g&������Z�=M�sŸf����#6[uX��"�Ǌ����TN� �h�)�U�Lk����q���_6�(�tz=Ii!P�Ը�&�4h\h5���������yE��կ���ٽ�{X�#�Mw��]idb7o�Z�K3��D2�y��U*:E4Ҳ	(Qjw��S7�E?�[3�c0z$F��;Aù�I�pbA�[q�]����fĽk��v���/LZ�7g��X���/��S#���D2�.�s+c��'+؇��Y;�D��[+8��#����pYR�i8J�AiȮp��B���w��1�r/�U�	^�`��o\�����V��'���S�S���'k��T��pp�o����.�:X�N������O@���?$}�<�����.R��a�w[5<���n���jT:ܭj��Vs	�3=:�w?�� cI 6��	�Vo"&u���k��'�Z�C���]�����kv��wx��^��D�s��rп&�?Z�<z�-o�Eɠ��I�� �e����DU�+^CJ�V�f�f�&�G�)�L��#�w�������4u!䥋n=܁��Z䊍GX���x��<)a_�5~��`
��M�B�d�)lf�j#�y�����]n!��F��,OS8	ub�,��ﯚg���}�H�R
��TD�	]^�%���MO���R(������cp� J�u��-�m�p*��=L-H9y�Z(-[�����O�����N��&�*�-�e�:Je�Ё�fh��ᅍ��|��ӕ�0S�3��:�G�
�If޽b�%�0�:�Es̜6ŀvDW��(m'�vw�k+��R��Q���R�i0at_��	�)ԅ�)� �2�/�+�ҿ�_�&+Bc���-�U��E���C]R׿O����
	�X5G���Y�\K�
�iJ��G�l�@0JhT֭+Bo�ZU&��,�BU�#螙��e�p&8� �z����MV��诋]dں�QG����\��F}�:k��.a��]
�8�;��%�H�"�/!q�K�
R�FȷK�$�4��h  Ӗj����L↶��u�����YmD��RT����ۈ�k��~ܗ�T�|��d4�y��Xk�Y���3K���.��
��o+�F��5�%�hw�	s�ŻY&3�#��F��u5�tج_}&G�Up<��r%7 h�D���I8�P[m�@~6F�d{��4�g�Gj0٢��Bt<x�kN�C.o���hL���Vl:���f���P�#Fb��30rvv*�|S����ݰ6���0�n�4=��sfNDET�T:hq��qbA�|�Ƹ[	��i\p��(�^こ��-� u�z�莬t{�s�V&�'�QU�㺯��h��������9�Ɇ	6�ŝ~
*��c�T���:�#h�@�u��4/Y� �q��z�]�`�}yIߋ��M=]��m�H�0���ۙc���m�i�;�9��s��]�C+ *!�5���8@u;"�J�y%�ۓ����|�pk�Q2��nL��~9�u�:4�;h�_Տ�t�[i\�앆 a��'�࣊%�	^ �÷�����5&�(u"�5�x=WR�$���ԙe�G�#4a�j��~�Z$%V7��j_7rP����Z".%��y_o�km�"������Sh3���0p�{
���lMǎ�m���#:Ň�a�_���-�4c���eG�f��ts�<��x��rǃ��z̄��C���J%�00��wK�ml�BP�O��ֆ��z��R���f��?J�KP�C��XnQNN�kQ��m���x�`1���Uqt ��ŷ��g� Y�3|�,ac/ U��P�x�3
���4A�9��z���.�g�vn)A�����y#Mק���������a�X�&�$Iz" h�LS����`*2'���qR}WHLL"�|����eڙ	tK���k�q,p�����-���#�ˏ���n�2Y��p �,|�.̱��"�=��pJh=**��͖�yYN�)�]~u'J�m�(.c�B�D�����#�b�}H��Gh
�b���^n�]�𶣡�D�r~���Le/֗�Wǰ�}���9ړ��_�{OO4�'��d�����1Q�����Zh��8���"A9i_&+��&���2�W'T,7��#G��z��/7U�ٗ��!­㯨I'���?�vQ�v�����F|�[�=���X���	����i��"���K��2��,��Ar��=�;��џ%'A-.Q�ǽ�Oր�F�������jpK`&���[g��F�N�Ak(���])�nﲑNKZ�<�n.0�`��t��f!��S�����9�� D�d����5��Q�3�K[e���f��7\\�/p�U���6�v�K���\��HwN��qWSezI�W�N�P2����1+4�9ul�^�� i7v=�X�o����rĕ��V��}��f��ȧۥ�}�������U�*|*�W��i�m����?�ى n��t�[Y�2Z��]�J'j�W0��z�0�0���=L��0����Q�r:�w��vn`!5_h�bq���>J*��=*%�e���j�0�lb7� �
�W����%&�|�^��J-��H���B8T�"��P������l�zC!L8.�$�D�O�U�7���A��5~��X<	�o�`k@�=�QL�'N�t*)�s����r�c��HF@�X,��!��=9 �G~���YSCtMX�^2��U��U�Soy�T��Y�&����[$΢��q���>F[�ҝD�T�4O��4r��/�|au��� �^���ñ�$�c���UtLf��mQ�D���Ȕ�HU?U@�/FF�<-[�n��&z�cSgS�k����������y�+�4�!����W.f#�7遼��b���V,��)�P��n�jp���bD�,�Y�4���/x> ޽�'Z}�`����O
��c�NF���qL�H .���?��-����n�j�C)�<��OC^�_�?l�q1�ugd�R�,��8�a� �t��2Y0��#���|2g��]�T�p��2S�˗��K
�T����t<�r1=�d���S/J�#���9�;{�Q��[�� �ȕmۨ4q�LpH�v �>�,�ڈ��������I�@T�>#,t��
�<a�:	��rS�?�N�&�O���d��%�����*��R*��w��$�.Z�G���#�Q,�Ke]@��Eޞ�՜4p�O���;�� [�߸�ڜ�jyړ��OT��a�G+;�I��O�gH�22�p2��Վ�,M{V�҃mF�F�֭��t��@�0mQQ��,t�*��3��jJ��B\�L��M}/�)*2*=�g�]�拷�0$�����FI��ι�r�/r��`�a����Ç8����lW���\��.3uFu���#��a�$)�2E�n��[<K_��K��O��Ɖ�"_����%�X�vN���z2EL.�PO����LvZ�F�>�
� �@���t^E쮵%͑l2{��N��,�Mn�d�߼�ҟKZȀ�(R�'9Nr
&�|�� ��͎Uf��nZM�.1<u�ѓ�,���M�t"Z:�=���C��M�W5H��d��En{��λ����N�M׼��TY�yT7>s�'�x8���'�eۛ6�ؓG��<�2��v��."�>Y~�0����7|�98��%�T�s9t4��unZ�[	�$��]������`{5��x�@���ft'�>P�����{���e��@��t<�bB�
$�%�=��*�n§�[����N�[����{��́������S�Wk�^2�К�G��${�P����[���z���FXԄR����ɢ������}4\�"�w�m@pR�v����ayZFJ����xH��J�{q)�ׂ�C��-�c��FN<��<�bb�9����7Ol.T��/#x�cf�\'����6�:�vV�ւ��}jU�s�9(��Of��F6���M8FY�Lr�W9���F�n�*ۺ���<���=�H㦎��'B�p8˂➋��c��x����O�$Wuո���'z�,*�`l�#��b9:+�j� �h�Qo-?��6S8���M�[����<8А:�)���6Z%���s���,���������)e�P�?����BA��b��?LCk���0�ZH^~�ۢ�gWg���{�"�{�ǧ^��A�0����f���a������>�SQ?�Պ>�+���HH0w��stRR_�H�2�M�*��|�;�Q�p��{*/#�3����I��<���n��5�,��ƙ}�$�@9���P���\n��?��8�T �d�u�Ł�׬ɳQϑ�X���Q���\;��J��FC�w�)*ύc�����'�m]M�&t1�m[1]�<?}Cay`�?��z���K���/��"hd��=��H��b���a��g4��۹s6s�26��C�5�{��R�K��Z����.�����tqdѱV�Q�FۤZ���<���j����$�e׮�'j8 �L�햜��XG��dݷ�hAt�@��yPs��_�&"���WC��b� ����Q�@����j�$ώ��Q�?�|m�G�#�@�ӵ�tM&2��yb����� /,yB�Q�E�a
�N��udٌ�p��_+`�k�_Y��Iۖ�*����10�A[�Uĳ�� t�
��,hC}��|�\�R��2X�����ϱ�M%p5KLQ�B/f\��ጺ��}W��H[R`��w�ħW�
r�2��Q"	~�p������׃�D����<?�W����#|��7(fTC���}���
����wVn��z�>#-go��\&���Xf��F;�BZ�.�-A�����ƕF5u��k��;frh����ML�Ϙ�%P4&a�ʿ�--�x����.\Q����{@��kD-��l��%����j0	`�8w���"���7����� X�x�y�oү�yQ4�!hX׍�����mX��E���kN�� H�3hA��0����Wc�R�ǜ)MR E�b�iގ��\�Z�l�%(�>����8�>|�!^\��W;K�'m�`x��ظ�e�k�ns�4VӴ���J�d-tcTa�Z��bqƯW����{<Gb` �����]ے�:�����Ɔ֍�9�Ya�F9!�D�,W4����&�E�c���l�g!BE0C��h�A���.ս�a�U�,����p�9Ȥ( �������[尅���|��x�p&�Rv�������% ���M��p��� oW�9lX����Ŧ]Jv!��U.�(�r]X�S�5A�~t���;J�'����N��� ����lQ�s����|�X�j9>���x�����V_�^���b���S�X���3Y������mx:���T����S����[���ć)X��m�	d��z��-��������dȗ7�<����s�bo}�|#QJ|\-���A��^�
��q�&��H��=��͒6X��,0�o̞�8Ӵ�>� ��0B$�����v�,�'7U�e��銷��PX�k��jx������t�(�7I%���$�s3}�|��a^i?u
�`j�
*Z�׻��qJ�s�03��<ː����o$���1c�h�w�$|���X5��W:P��F_?����偟��`��-Sn`��`e9x&G����&տ�خ��A:��!]Y$����Ca��}��-��#f���wi��PC�p��<E#�φ-NصbM^�qj'g�$3�:�S�л���M�Y<z�߸�QƂ/�q���oN�C����c����������<JU���1V�L7u�^M項�����Oy�t�%1�)r�+:�"�% ��K���Dcw�Ʃ>�>��R�w-B�\�O�D�Z���A*�/T���*O��<HIԋ�2�Ͻ]�c0�Ĕ: �����i�xU��c ��se���d�]J�����ts��B�xi��{�r��$����N׆	;�0�vI������Q�-�n�K�O��C��hq�R��W�l����Ha>B���\Z�_�4M-���0��}+Q�����@J������0r����h�de�X	��J�v�����UZi𹏂��t@@P��St�
�w�&���+��_�]UTP�+� �A�L�@\�޺C2J���b�]���0�d�eU�}Z:ϟ>Tu0��5�Vz,�0��2cP"��k����[lH.0�rr@�a��^��4�<g�(��}D�R���95����&rR�>��_f�d�`�Cw/��-l���]g����g��w1��=�B`Bò~�o��@6_#�$U�ģ�N�d����9dwѽ��Ʌ3��m%*T�c�,j��ީ���®+��[U�8l�s2��������x[l݌�N�����j�0K���4u�f��g{�u0|��PvK"a���27~��g(��u�"�|���7��L�|��g�#|��P��3����Q�"WQB�ݲ�h�	�K����JbP��`÷:���Y/<���l�H՘y5B��
l�e\[�����ȍ1�;�=Q��D��!ױ�+�:����;�Ӗ�D/�q�R�O���eM��� �BKS.��)r_x��X��`��,n+���8� �>�S%�&oE�moXY��Dk�Gsx���4�\N%�T�*!�R_`hb��BA���fHS�R�JLw>�z|ք�ɡ#�̦Z��\�_�����
h����3I!�T=����;��M���&Zv0I��a�C�?��)�1��I���kV�Ӄ+���ë��!˗�(���( �.�y}��X�'������P�r�����@"����ntLUr�5��퟿�S�&y���gudA�j�:g�w"�h��n�Q������3�\���"�{�Di�����Xhk�����oxÎ��N{1]h�a�;i]�ޓcJS�-�?''�T=�I��m��4���t�'�t�5k�+#�Q,�Lu��,9�z9�5�{�ܹ=�%�:�,V%*`v�A�|����C{TgMt`�'�m`���܉0"��)�p���?JJ��Buy��Hl������S�#ߝM�cvO�@�r�t�CU5��"������MÎx؟f�(�w���8�\,��Z�X��@�5rw���ޣo�����6H�2�<����8�@�����Ssc�3ج@nlq)Y0�N�)��naO�@\V��ΰ�y.�瘼x����U��@��]�2v!����W�Wb�⦊�lM���ez��8���-x����/�$�װ궂�4�}��>;x�k�ڧ�����!�a�<5br�WIHM~!�xR�|���z��&���ݶk�L\��m�$������N�2�wM*]hb.p��=@�wU�8;I�{�ȒWЏN-��Ʒ\��4�ۋS��!K8 $F���d���))�lk���Tqr ��oDQ��$�>��� D{e�K�Lt�[�(t�������f��'����*<��ܳhn��a��'�!tA@}~g�
P�H�ڊ>Ao�pAY�
�'���!�e��%�r�T��0̓��!*���/���5�0�\��1D5�+��',�ܠϻ
 7�a�)ն�#������X�$Gv{lf�>a���A�WYz��;� |M#�����5{=�К�ݐ�F�W -�k�B�]�g��r�@�zN���Q��~���`꺉"�y��62ێ�f�)�>�ޯ�L�[��s�8A�x�������I��zf2>}X=LGk�R��`������T%���Kz�kMNP�Hf��3��Q �(6XVƻZ���5�/�̇Q-��nQ��ωG�.��>��r���Bpx����K�9v��(z����؟��KZym�>����=�Gh
ϙR^�?c_���4�T�Z�qOۃg���:����&���r�e o��*�7e��j���Dv2�{=�?aC(B
&�����Q/Yr���9u�����Aq����@���>�%�TV�:����'� �Z��$Wê4W�2=�?
����B������\�i>��� e�3Χ�l�#d�c�� j���8v�k��X���ay��7�U���$����qՙ����Ϸq���#�
|�"R	��`� �~s��E';��m��+\�"�=�^�-e����n�hg��y�4K���G��e�F�m�@~�O����2�ˣSLS2���V?�`E�P��E#�^�kA�5����I�;r!,)�����B�F��.7��м���g��+{��
fu�I���㫽�;�/?�����Ͻ��� ߝmeT�9��٘a_��hT��Z?�8{V�Wؙ�j����!�C)�:��oЗv�8����nEH8o�|&D��z�wR ���1��ʼ�������(:�J���h�tͺF�K����-8F̥��N[�<�w�^���~V}��v�@�_�OJ���z��#���.�dJ2y���$�C_�����+��S�R��H\��%%�bJ��ɖ�cy��[��M��T��~=٪#�E#�`�t}�Q�T��Jn�W�j��j����EMXPl:�G�)��Tޣ'��Hݣ�o�<)3�N�!��f?�O�=ɇڂ(wi�)������x����~��	�����[�E�v^�$���.O 5ƈ�?!+�H���8�)Ճ��s�*������rks
*g^�NW�]*U�1�*��?xj�4���#6���SJ���)��d��z�̩L��>4Xq����35=9��v�y`����u>�2њ�Q<��&D����%
�������c��-�{�����Ұ��w����X
d�m��%��d��^ꎑ�E��A�Ƕ��-v"��p�r�����U	iz�(��p>Vg>�O����kIC��,��(�!���q�u����ܘ�'S�*�4�;����$*-N�N�h���1V�H��~��{�g�������@^�_�8�秱�B4�t��t�l�d����E��3jZی5y���3`!��ٯNF��)|MT��!�E%1]��R�q�Ȋ�P�e� ��&w7!�g�:�M�Z��j6*�zruMhW��}^#�[�SM���p��d��<��5c�*�6޶>�� D��w�rR<�8��!�#ض���ʶW<wC�Lw��<(��������Ĺ)��%��Û\���$����ʵ�bq����b��_�#�^�c�n>�{����|�U�0́��u���6��U)۰Ǯ+�R�L�GuԻ8����Ul�/�#��8��������Ѳ�T%���%)P��a��vCd+���S0z:��]3H�1����W�\(!��Bg��QIÅ-�d�\�aAD��	�uj� 3��9�S��l,{8x�Q|M��ƈ�E@��U-�LR(�7%Sk�����b��M�ϣ����� zD竩Z>jOO�e�U�T�cMJq�ЎXf�"�Ay���b��iSt"ZO�&����st z�_�����<��f�2��j8bt]*	���5K��^6�X��6�G��Da�c1��m��<F^v �����J|W:��-v	7ׄȞ�kd9n��O-m��I������ ��� ?�a?e�}rRZ�B�P]ޙ��~҄�s���0���v���� |�z$�С��x1�6�HKHp�l���mi�ͥo��ˏɨ���/���yZ!D��[0,/@�v��E(��j�H�Z�S-Ԍ�I��/ z��)87��>�cz �+|?�@G�%��Wq],�?ݮ{ �쩉5�X�U�[`hH���r/Vl��H��P.7W�\"O�ˢ�� tb2Ԃ3�b҄s0DX�oTC���Nٿ�y#8���߱�Q�M���u��oZ�0oXT$jɱ�g�oN��a�D�Rȗ�� 	I�#�U��u!�;��@UeE��Q���M�Ԗ��,Ҕ��T
��K�J�q ,1F@���}�,םC��ޏ���k���l}�_�E���oݬ>�D�=��#
<�<�hoa�.�փ�[]�`�����ҍ�"�]�p0���q*�{.ز�Ol7�Υ�sߔ���9�~���aMVN,��.]��!Z�<G/�q�-�����K��
��s@�h�*�b��~*FaR&��� �ܞ�F���0�����)�2f�7��&�{Md�D�-'�(�}c�:=JQ���^�����c�k��Z�?	j,UN�����(*����1�sj�̅��Q�^��BAB��e�}��U���\�{�3I��xM�1�"Z��I�����v/G�z'mf�������W�Z�JO&3f�Q�k��4�#	^Q��t��=!/^e������Ș
ϥn&��١v�_ܾF�\X-&/��P�x���	����J��$
,�F'��� t��e6d"{ZJ����9f���40/�ǧM����a�����hG�_z��W9R�[s�,�3({��6�� |V@Բϵc�LF�|�:�}�M0Zy�R�c9��@/�X��^��>,���4X�\�!C����x�OV�"�g���jZ��O<ۺS\9LRK�N�Ԓ�p�]0A��T�}(k�%Z4��r'�-ZO1�[��O��T >�ݢ� �A2b��Fߒ�����$�s�10i��v��ܯ-����+���Z�磶�}x
p5�]���y���{+��P�[����ϦZ����S1���.�?r��h�×T�A����Zo#c�Or̶�歬�q@U����[��K�|���Y�����	 ��]�7�$%z��;�����<���@�z��n�	�u⠿��[�Z|�8яKk8ɧ��}�3�g�)���hrގ�v�����2)|�v�'u�4�Ze1�@H^�o�ޢ e��g{�~��>�W���6�HL.��x�Y>�������v�b���	 ��cMO`�D��&JR��}���&r8�!�&��I�fg\	}�	��5���6�K�&I����ٷ4��ߍ����;S�����ag�L��X�CZicӰs���@��U�S<3�S�e��K�^ӯ!Q{Ky�,$f:�ɾ#�oW���B����}�DC����ݕuY3�M
Q6j�1ړ;���ܥ0<T��*tO���`���|"���$�~i6�����\31�C��1ͯ�����~��-�a̶�B�z-�%qr4��13Ξ����=�O���Hdr��ZD��H������GXlW�y$�U�q!_��`_M$�M����(�
mk���3�Ta�rbM�?�&9�ˇ�2�=
����`��SI?�k���X�|'��?~�e���X�i�\"֡��� ��J��-%���1����[ɠ8w�*�5�~��Wϒ���lf��b��x���h�|Yٚ�.��?V���
u�����>bs��b�m����w�c�j�����x"��	i�l��#\�2��׺£��8}p�Z�?�H��l���&�D��5�(��:��̂S\�p"
��ׅM>��b4�������eg�� �sx�ȞڇG�0��J�ѐ"(t���Y�o�j�1@�HΘ!W�{?� _����%Gߝ2��[y<��L�cB�8�%�e������o��>�B�%;P��=-zE��i_�W
ps`
t�z�[U�{�=-��W^b����8�`���-���a�/���,Au�E�u���VAB��$�y*���¿��w6�����A*#�_�f�E#ꠟ���� ����V�h
��]����?'*�-�Ο�1l�lt�ؒ_��?��}��n����q��ҩ�m��u���ƭ�(�S�B��;|��!�
^�_�a�i�ˌ�E�; +Q�'^1�������Џ�!�h>������$@B��� +��+�z��A��(��&>a'!D�uǑ���i���[�I@<q?�F���WP�?5�I����0�eo�_�A=e�b���P��@n��<[��$撡���uq�޸.\z�I4�uFͬ�`�v�dE9�	8%J���z��xBnJus�ռ޽�����4�S]����;�ֱ����������r=��O?�~�t��Fu��t��,�$^�Գ4�0�\n�	~(l@*�Z�t��W'�Z4tF
�:e8O�t]��&g	m����l�����p��8�H�^��PZ����s�`�lj}��m��К#h���b�����KA�zpuY"�R� ����67��I����S1�]Z ���)�sz��8zﾊ�4j�b�����[;�yW�b!�&݄�<}N(khy��/\,��]*�����5��m�J��R,Ǌ�������f�-i��
�Q���}t��-��& ��[�܈�OD��8�*,�;���k����Y	�
nc���%�?������?���sEX�����are���k@%zef�j���|]V"Wd�b[3qi�#W�Ö<%og���Ԥ~�������+��v�u��Rng��V���x�0���:�*��}�t�Q6=� I��S�FD��7�R���h��Elz
:�Z�1�Y�%$o+�
�"Sz+�Ÿ��7����k�@��X~؁�-������F�
V���b����"��������/sdF�N���/����m�,��ūj�?��;��[����W��ú�QG8�1�K��F���˗K<��C���JH����Tй��"Oj<�rrO�3�H�'Id[H��9�WeRs6WB�Q��%Igg;��X��]s��V��[Ǖ���ꂬ�5��J��cN��'�]z��dX��&HO���X�;7�i���GJ�������Մ�Е"~9-������~�ٻ�l��z�J��+�!l�.7-�[���XQ���b���'h�'�r�AѫK#ˊ��H���lA�� �|Pnl��T=��=�9����&���G�:r�U����gwL�/w�R��P������d�m�Ae�^��q�M�N+�Q�4���p�y2wkQ[��X�w4	�&؅iC�D���ȓ����~���\�ݭx@�8�p�Lۗ�.�<�ѬI��S|��9nr���D�x�L���J%��.��1�Z����Y�>k�����P�UA�3����Bܹ�$���dFg�5�Y�m~8)8����>���;,bl�I��uf�0�p�b���yEQFN*�0���M�qKn��J�?�
:m��4�=}=�p�1�1 �S�f!�	d-��?��oA�o)�]Ij�?o����'�_Z��Xeʱ�)J����AטY�I�wlt�e4s�Λ��g2����.����>v����S��B���
���WO�V�
��B� =S�V1��o	�q'�Ռv7��9`�� �
�ļe�d%�ɮ|�J����'����J�	4����D���e�r���hS�n75vpt�0�kX���\�S�oZ�7���Q�Y�$�ތ�`o��/���^L-���O�@�u��s�,�oX��U;�ē���r����7�f^"R�H5������d����D2Ɲ-DI�2#�-p5�H���UQ�X��=k ۱�HxX��"V��/�~�x?Xt�CM;!j�fXa1Ȇ_2�>��/�!����N!�%�)�r�@g��Y�H�63L�B*H�-���>�M�	fV5<�[�"y���kJ���o�w(U9���9� �X�|�&�	|:�X��pM�sç�m��{ٲ�y��l�����u��#��m�Jz�����=x��w�zl�EN�����s��{&��\��{���|V��*o�M7X��MNz���l�48�2��T��|e[O�k(@��%m.�m�YE"�ǆ�Q=��z�4���Ҽq�o�7q�*!p����i��$���c[��CS,6��7�(M��-���Q͠q+��[��c���#'w��K��n"B*��QG���"�S���O`Z;_Pp�P�����iY�Q-p���RbỄʔ��)>9n������t��ي�M��U/��*@&�'MJ
\�p�D�Js�W�#W����ǂ�E�U?wj\��1-�<�w:!��e�Nڙ�-%&���L�zk/f]up��v�AX���p��>\Y�u����_�!����\���m)"4�o��N��]��>�;��i�i��k�\(������A�ŀ�D�.�V9&� 7�>������`.��'�r�hX"r�j�3�t"���ezl?F�h_3��r���
E����I&�0s~�+�/���i�Z�43������3c�}��(��RX�kI!��OC��C 0A�I}9}Oe)���\�����i �9��Ym�fo�I^(	'V����Mf�4а�+[��^jS�7"
ㄦ"���(������?9q�N�����dtD����6�_�/� p~�z8>�c�#	�k�j^�wwG
=�|�֖K�{�}��SR�a����̇!�4���R����`:�N��,�i_��z�2(�q�Ē=Q��<��3�"����@��Ԅ+�������K���������]ʷx!��u��p*+�
��>�n���$7�">�/��3��	�ƞ��	l���~u�ZS����ু̝w�K7� �.!ج���!��۬��w����,GC6s߲�t���wL�T<�<���D�:�b���?ȫߵ��â��au�bB[ ��?
$�~��EGUŨ�$�66}|��F�40���4%a�{ы~��x��v���'��V�|Y����i.Y�ߏ��"�c�O�����s�y���/� �Gs?wM���W�:�X?^('�U��������!_�g� >���/�'�0�v���B���Y��l&e�7�T�Gt�F�4ۜ����~яd�j�ؽ�ȩ�C�ň.����`�_�~eh�G�)鸇��&mg�݈X��ۂ� qF8"=��JT�����q�V�|&�J���0��M=˭��|ZUflt��Q�����l���"�,cP�b����VP��G�$-鈃\���8�}�")�Ls-�Y�"ԣz�D�k�w�A(�C�c�B�~(&þXj$��f�겆�	�A��uz7$=�f���*心��d��o[z�\�>%;#0��ه�v%��@	y�\����q�*ơB�V�C�A_Xh�cW?:*HEGIzR�xSAس=�g�BO���d�N:��8v�'��{��v3�M)y�=[
���&sNE��dg�׉󋓯4�Vgŉ�=!� ^H+�W@=d��C#��W�)��)�NoB�ߜ��(���_
��GC�&~vV��Q�pXI��휪�'�8%�M�P6�/��X	XU���o|�^��J����/v�y��z/��˷r).`{kxv�	"#�c�WH�p�<2,���������Z �ˉ�G;��Z�"^O�T��Y�B����1��ջ0ڽ*�g�5v8?�QY�{1ڂ��<��@fu ��L%��̕�lHmdd�y_���ų�a'
U�/_Ky�r�t_+�ѻ��$������lg�L����25qnS��qᇩ?�}�:�����`7GP��}�{�s��l�V�ϟݣE\�&a����}��v��i5�S��NԨ�!�ĭ�&���BHxS�5�5���*�"!�ƧڼHU������� 0���Q�z�}o��{��xeuc�����m'X�heP��&4R�;^Ȓ�g�$O9���w�9�ߊX�������w"z�$τ���Fʿ�4@ߘ�F6���ȭ�Y��zdW�N�r�_�=�LB���;k3RM���G�����jT�A��9}�VX������X��4�u�T]�h-@����j!���'�l��P�I�{b�S�		*�Bռ ͔�>q�L^/I�?̿�/s ��=d�%]��l�F���!��1OS��_����#ݮ� Nb֑ }#|��5��[���8�q­�Z�D�ӟ�[�M
Tc�-3��5u���	;%U�)%m/W������P.��Z� Y���h�:ڵ����GG�oɖ<,��Ɲ�]-�gy4���q�.fj���v��S�d`�+�׺����t����|��]5a�l�~~e��hkTFo{ZT�!�p����Q�3�Ms����	�Yd)AJMmo�σ$�K���V�s�Q�{�쐙�"�W_a��v/ �A�x�6�A����g[%$��Z%]`���87Xu2]0{�p`��q���V��HFq��6�C!�N�t@ "n�Mn��yI����"�~�*���!������Ƃ/y���\R�^	%��������T�|y<�߇A�̮��m����U�-h��Ǯ�9tvJ�I�AO���w+��e�ᛑI��.�k�"�cKߚ���1�Mԕ0��-�*��^�	W��%z�NÄ��΅}�L� LH����&�5�0�N-x	u�S5mu*u�o��K�yV�[n� m3�\1
�5LG��~?
��o۽�M�w��#Q�V�[��6�j3N��e�P-Ed�D"��*[���CЋ��{ɧ9ѳ��؅x=7�IkY-p�R�MV�2���O_� ��W�!r�S5�w�:�	D@��zb&u�B�P&K@ר>+t`.��R|�`��Fw'������?5�a׭��WsMz���#���iI:�P���[[IE�>u?/z+�tݚ�N"o�*�d���3z&W��t�M�G��C��M����������-�%�\Y�E����nKCO}^9�)f	�& ��
�@�ky���(>����w�RǺ,P)ٲ���	��H@�G����r����v1�W�*}�\֤Oa��O�g�'��y�`��-�A����(.t4��Tb�oSu&��e��r���h��bR��E?-���c�l%�2K�٩D ߻��$}�[�R������<�<߅,^�N�DhS8矹*��E���̾��k\җ_O85Q��ˏ�V��M#\"�N�|Ou7����%ɑ���+�=�c�c�>��,�0>|��r�bR�պ#�ʛB3�=�K�I�ʑ���x�߅���u$���N5�ʎx/t�q)�Z�����<ʟw4`s��~6�G5%�d�#q�\�F���E��+$r�dE�ƃ�O�����t��=O��jX`��zQK�}2,�G,ɖFx~z���GSF����:�m�XL������ˎ�~�@	g�!W�Fa��c
Ō� xM����ATZl�0�f,��I~A�AX���c�(Z�tu�dTo�+,�:�	�Px_��s 1�0����+W��n�}����ئ��}x��j�3g��h�CC�/�"83G�`����}�b�F�l��(� ��KޜOR�6,�邞��Tů>~\-�7t�s�:�6Fp��&��@���p�� ��r�B��*גoO@��ǧ��J��&�V���ӂ��	��7qn�hS�f��]�>�Hl�P�6.�|:{�qQQ�J��iFI���t�5g���'�=���Y��(ȭ��g�� �o����.��<dzUh�32'�jrxG��$��E	�*Z��c��+�ڣ{
�����G~�b�u��1|5h�eC�V�=Q��t~ 2�%I�ܥ�`%wX��D��r� 0�����*�
+���l�Al�%�J+��I���Z�	c�XM'��S�M9�������f�u��s�Hl
W!�Hk=`��3�+�k������� ���	I"c���\����C����?�� ���'y|R�&�bU��jt:��U���/6�c��*�]���$�p�����gG�3q!zZ�D����r�E!2��&�'�ɮ�,���9�enx�%�xe�^D��#q��"��z�g�������]./֜ ����!ԣ���XsK:�0I�,<��)Es�����I���;�O��V�,���a!Lo}PE�i*�N*��?a(���+H����A_�- ��2,�����0��1�k���~
��o6g�ѭ��6nI��tj��Ԗ�jR�[ԸG�F��v�Bh���BM���Yr������S����F�;����%��v'�����&��C0��o.n�m;� ���߱L,F�tJ��e���_t0+7J��3@�++�ٚZ�Mk�]�����1g� �}���:�ZN�m�N5�<��r�h[�nx[W���3+�jq�v!��L�3n��Hv��.k��՚qk�2�h��
�����������X�a�*��H�G�p�풵��������zǛ#�i��ȋ���ฤX	zX�p~��i�_bd@�LtvF�4�c��������S�]�!vI��>�f������� 7Zx��w�Sk��3�h��KX�i"�
�"��Q��Z������?��ѡ������$�|SL�p��9�?���A9*v�F��U-�c�Y:���ݟhh�nm��yrz�G����\�3h纂˼�uƞ[�E����`��Y�l	}a������{K�<�����l'�J�L�9x��S�SB�6�vV��|�8莊�[�H�����_���R��%$�iVh뒍��#d��] ���J�H8���NM��:��ϻ]<�}� d��t���4��Y�37�%�~��f")v�&���[^�į/�GW��9��J��@�k!W�an����)�"�������� E��j:���o�$�>{��%�0�����5s��W�Ϡ���՜�w�-�K��Xp��-B�y�G��T
�y�N�O���r;ij�v�WN��(_�x��&����MA���TR��'R�+\�7C�#�m'� A��<�Ɔ_6�_X����Rvp�;����z����D�W�k���9�����n%�N���$怼����؈�����F����t���V���P�Y�Awd3�F�(�!���Z5�S�Y��������������l�!���0�-4�5�%�W�P��l�cw��f�؍��>����j��*6��X�����􂵥=�z�s���������+%2�IԀ#Hx�y��'��`~\aM�dt�ޕ����.*�)]�f��Ժ�~�ei��j��_&>�E����>@T+K0u3�8�TO�x�uY�qP����$�ǽ��8�F���c_SO��oQ��D	^��2iگE�����X�2��N�:�Ӧ�*�)T4���@����]1OF<SY������[�Դ�e�O��^�	����M���j6�����/}mxEҞB{�����H0��4�nP1�ICH�j;��F�i{P�^]�7{����/���j�CW{�Vx�ĀV�2�E'�Ew���r��gB���G��R��M�erUo0DG���ςB�jlTW�n��?)@��͌�ء�������h^D��ӛ.{J�{b��	��+@�u�}�;#�Z�s�kR�X
0�w1�ínl�uj*���]�Mh�t㲀�\�9;H���{K�>*�B�g��l���jң���,o{{�j�K2�7�O��L6���/�x^��D��,�����A���X
�����%nEdP����*��>U��6�j���G�ft�wFJ�?)x-E/��'�:��.�޴�I��T5�k�	��("�P���
��jd�9P-Ƙ0������	 =�� ޯ/�4��%������P���,�8��2[�"[�zw��/!���	���A��� KA���]AG�׶�l�#<z��y�Ł����:cl���AYk?����ւ ��W���g2m������4X1�XZ}Y�7)�
�n�FU���'��sxLϑm�6��� ���$�q�{�t��|���@�n��$���-gNz���;��<�`_AS�"ޅ���yĮ���vجi���`XR/��\޶u~� ������„�D�]G]A�yp��=�Y�G)��&~J�HzV�/k)F�1r�l�hv���������<�d���V*\`;j�8�TH�b׸F�Z?�B��E}�����:Y;�̺F�,, V��.D�$�=g��/<g�"��V�_CJ�����f'��v�����ZMF�
h�&-��z*�;=�.giq8ٖ�3� s��,����+9�r����ڠ��a�.�s��jj�P�9��Һc+o-h�d��%\�����f��VQN�6e�1�>P��M)G{6&�������h�,��3X���˂���a,ai���v9iW���sJvBߝ�|��n�i��lV�d�4~Q{}���d�fq��T$��o#QD`k���=l��>�`�@+niݰ b�W:ͨX�������v��+A>����������-Cԩ3%O���oֳc�X�u(ICt�9�L���B$^��\<)���o<��{�uJ]���l��<}%7�����p����l�
�Z��,�E9�����&.!���\�R^��@�����0��
`��g���y�la�,�� �w�.�I4w�o{��� ���Y�y�i�K��g9�jF� ��o�����vV�ٶ�JB��;g��S�T�MR���,�_�Ms�j�B>�q�k}�	�q���z�(y�K�C���_)02��ց`�%���N9GN^���kL�fSd&�R��� E���πk>�y~�A��t��3�62�(�6y����t]�� {�ǘtVa} �d� i����4��A�@?7%���D�k�Rt3����1�8�>(��� `^6��;
�r4]]( �r;����#����OTA?��E���O�'�"��ǹr�]���Y�0��TZa�y^�2��� _;b|±`-^)����?ʵL���Y��夰�fJ�.A>.9գc��Zo��=��b8-�:�Y��I�w�T��n�|Y]�懎�
|"Y=�8w �5�ƒ>�K��t��j�^Y�l�(�$����.(�z��;f��Jj���p|�UW���ұ����DXi�:"���9���7�yϪR���������  vW�X-�d!��\s`�E��e���������a�̖o�fI��������t'@u4ke��^(�M�l)�`�$�?�<�S�
��Ʈ/?�v&�s�9A���O�R1�9�i��Xl� \�4�yQ��� �Ⱥ%FY��ZX|y��NK�(�����Ѕ	��G��JÇ��j�\�]���������Z*���`h���X,:$�K1MY����ɧxE�@fl�f�4R�_��������[�}���ːTY�+��4���l����ܘL�����}x�<�c,�0B4�P����"�)�w�X��׃�Y�Bma�~��[����ɥѽ�`'GN[+)�'��']�3�q�>�X	5�k�3֨5�ZD�z�@-�bp$����	�C�e��6 n�@����޾��>��5�취A�)t�u��,���A=>c����	��/�D��`<�ʽݦw�MG��%D O�Ҫ-�H�����	@ oY��e��F~�fʛt�C���
�s��Q�I�g}Up�,{��f�B�]�tt�l.��8ƫ����&�u�C����+�_DcǕ v~q�`8��(:���l-=�v��L�{#t��x��0R�ճ=8߇)CېIC�1꣺)��G���L�д���"�9gBj|p.j(�E��NrG�):���+T/]�V��r��AĘ���ڛ��GR����sTzy&�� �'�Ό�0C��D-C"��-��K��ί��׵Aq!�@���R��?{>����1�L؜�G�7_�$lM��)��6���"߁R��C#�k�{B��W�{�����.�����1Ź�Y^�Ӷ<�F�ⶣ������ۯ�Y%�����/�zs�N�����s���8��M�I�B���;��"q����t����Ү8���jK�VT�4�~7�~G�d(���Q1����'u/���0G���D^-@��8r�!�徚��P��������ݨ@a|#`7X#-��.���u��.d��`\������z��K��R����*���]�H�Z�l�&����D>(>N(ҨPv���Oc�:�����rb��/�~�(d�~1�Z
��S
��J}�%<de�������$V��I�\%[%���:%�;���QU����=����\%����Y1s_nZ'5��?+N�I
ܭ��/��;�g,:�'��X�π��=Atϒ���ʝ�;��uI[�X�ȮO����qڰ,`o8�\GR����)I�筄�{ǻ�=�89����o��o��^җ��珅+S��'Yg7*��>ұ�S�5���Cn����k%� �!m;;W-`�XDK���;?�m��������j�q�����36��ڍ�HW��nC5��=��0;D�Xɨ\���140���Ԏr1=4�.#1m�(D�a��HL�<u���QҾ'�������װ��#���'Z ���HHg|������cj��m��9/�������O��Y'F�Q���`�:)��#�߰4�.E�g2ct���O��4 �i�34C������䵔��"����EQ�^�۽��5���r���m���**���S�?p@h=@K�#[��`�WG���$ Uk�X��OW���� IR�I��HQ`苙��D�,�J��/(��E�E����K�f� 3�2�� �2�.��(���<����+�O�Ѿ?��Ɏ��SL�'݂�*�aRO�嚗�T�i!�9�1R���A��(в��WB:�/��M-l�{M;MN<�%���A(?�Yr>ƭ���G���ء�)��Nt�c3M���i���~d��,k�cH�g�3���B[���@3ϲ��{<+&ǆ�o���A�%v=����L���ާt�������5���Nk��8���UX���pHC��38AI2ENK��/�2N��|����c����Yv�Tx��p7Q�5U�(��*ˀԕ�h1��hz�����v�oܣ��zK#`�f�K��}gN�wF)t���$$�uJ!�a���gI��7=�z��!>��^��l��@��%c�/.��?�ǣ��|5��j����"���W����t�`����\# �V�w|�;dZG�}iZ��V�&�+@J�_"}��D0�3G�XM�qޕX�RGVT���c�{M/��?֗I�y���'#J����Yn�4[�I��D'B`R�v���h�Rv6�S 3���6���|�3}f��8�}�n���F8(M��[��Y�2ո�W����ڳ�c��`������;�_5�?bQ�$�|ـ۫W��å8I{�D�C��3E9$o������d���3�z��j2��IB¾"+�h�u�[���%	�#�~kv���y^��.��x �1~U�ᦚ��5���7=����ػ�s[|2`
��r)�ڲ-�V48�QA����?���7=��[�y�6��C��O��gP��L&Kbʞ��@(V��_���6���to��>4>A/��raB�<�U[�����{��oU¾0ь���ń�C~Z�X8rWt{��!���WC�����ܒG�~9J��k����q�����{L�|Mn=,ٕ�uI:�i@@J���r�C5�,FOEm��I!�?x$�>'a*���������	��{J��6���q��֮O��j�s�`��$�}�.҃d����B^.c����o���g3�7'��1p�n4F3�AR��Z�K3��+>{C�!�c�����>�[������2Y?�p*��ߓl��׿�Hح��z-�=]�KY���~ ^��ꕡ�S��k����xg��aё�Bқ&B�X|k�X��$��i'���@��	9�$�����[:�WAݑt�3n���ro:���I�\+,� %a�]����f�v���{�K�y����oJ������tzpx�ۯQ������KL8��k����D�;��"����K���y��2����>ο;�ґ:��,2�&UL+�N�k+��hԮ��C�x�?Zb�@;��'C|-�T�1�������tw��#�c�H�?G|�Y2˱^�3+����wLZk�J���RZ��L:��oC<P"�&V��PP�D� ��������Ǝ���(�מ��c��[Ev�AB�Q���5��6b���7���1�uނ�?���Lc"g�f��Qr��g�2��ё&�c��ͫ���t��e]�A>�J��Q�@�O�+#]y�.��Bgc��^�/�"X�y��~��&��*�G6����������8%I�2�XyT5����~�F^E	����Q��Ô&e���p���p�n=-��X�ׯ�;�ڝب���� J�P����/_Ż�]�+��t�M$ejh�(�!�z� �u���D��~��wP�@$����2�\<l?&�����T�4:i������߹Q�(Hh�`]�ؕ�k���=��\��aph�肠�k/��`qS.���d����.���y�Z��������?"M_Kj^�T��<G���H�2�t��mMC�gA\�=�tSS��7k`af1�����<�f=:)o��L��w�"�)�B���l��a�
y~݆-�!�}��R�Q�gP�{��m�
�ۥUHb��}�yOz�J��ٹ��Rϊ6^{�VK���)9N/NY�~36��D��1lO�z��z���16�qH�)L��2x�>I�dY�'T�Q�M Xly<+��wIZ�C��u��j�U���ئK�zN�ԕ}�?��*R�åXA��VE��S_�P�#`�V�2#���O�P��HÁ	8�2�����|}�`!����������+��u����5͸a��#�xE6v)��K�t���� ��T�@�%吠�)���$`cx-^K�#�y��r�3A�z�Ei���E0��A���_՗��n����3*������1
j'�=鮈�7�5�L�)��4�ɯ2YtP(r��|��*F^>���4P�(��N�)�����X����z���9��)�Z����=!��e�n>�CF���>J�K��v�Q��&�������:�F��6��F,g��2	x8b� �t־���|�N,��:���E����ǹ���:���j����Q8F�b�W9��Oz�)Ϙ���[��4�䰉��	���0͘ˆh[����d)&�J���n�-2�2T\�:2�8G�>�yN�\��nͦTdЌK�M��XYX*��3h�xG���\B*��=1)�a���Ҹ�j�e/�7�WP�Ls*��Yd[���iK�Y���Ҹ��8�$eA���?�Oф�1���	�Cn�L �,���*�'���ƿ˯<q�!K�����C��-�`�)�/��u�\�0��qtG3.�H��G��R��
#�͝ru�.5�0t���z�)z���C˼䡉@L����.��׎{|/��j[�.X��ѱ���<>��&�(;��G �I��5`X��20�`��R�]��M��33Y*�v�ܓ	�!�?����	I��#��K@S�3m3�(�&��H�Z'����(�o"Sd{�Y<9�΋U����r��J	.컬���%+wX�y�}�a�I�Oc�u��_�g@\J�j�s)�#��(� �{�g�o����wv� �(R���zN1�0�Ů��`�yaI��s�G�8�&dHvmw�ߗ'�rVO�A�R �#whOO��\�]�_���?ZV�ta�c{t�"^A�"��c �{L�R�
SBX�b��]��h�hBt���meT)��Fnt�W��N.��׼"2)R�3U�����mf4��9mx,�?X���!ښč���g��+vP�I~�����]M��#�f�������Y�<���/�OwWAj/���EH�(ES�sb�pQ��{�PĎt�|�|�/mqq�x���~�ťkZ8��պ��PSH1��Ya��Gf��T���L��%'vM����y�"y�:�����޾��m���Mo���;����4��t����-��9Eb��m�fdZ�����v�XK�W��W4�F��ϵlZ}p`�#R|��.�o��w���?�0�v�����R��i����[q�I��s�W�" ʃt�v�{���2B��҂�*,��̦p�ֶߓv�,�>*���^�2L�RՑĚÑ� 6�0�BQ9�>MG����7V��:�t��|_)&\e�~���[��t��)�����P��%m��3�n$ch=p�̓;:me�痕�G�W�>l�B���-��o���`��C�����jo9�A��H�N�7�f����n�A���=��ޜjnT{:�y"��@r�uA���$��
�RKE�KۚFԍj�\��V6u��mA�1v�ԣNS<�{Bl��y����Q&��:n.�"���v��D��:H~:=m��{�QX�%�R�ʽ��:��]�hrwx�����?�{���%�
\���߽W��b���"�6�d��6��]��/�z^�3t4Y��Z���u���k�@H���2�u��Hz\��+w��J�o�* �����k+���8���2�go�}
�U5�2ޅ�x��r�Z��!��Q��1���\���*2���&����C�ႀ�ã�����`���Z����#��0��\�}>�x�E���n� �=���{!��n��N���p��3
��������~���#"do/c�W{��y~�>k��~	��[Ĩ������j���%]��$���p�VO��4q�u��K`Ѽ�ڜ6�E�oJo.V���HZ-� Õd�����2�%̠J����H;����{E�A�1	���"���U�Iu��'��]+#��4O�}�.����Y��rC����g]�D��z+��䑯��iGq������:�ǫ*�zD�%@HuǣY��S� �xN�]��/��.���%A��x�@ҁ��e� ht�ϴ5�߈���`�]��P����ZYq����Ji�Z��:5��}�f�u�ԟBQ4�C��.���V883�o�ٓ�|�hJ�T�Bw�4H`#{����l�&g���-9��Y@���=&��nk�qD �v��n� H7kOeIZ�a��Vaq����o!�O��'��G�X_/[Pb�7M���(*�n9d*޵��ʄHfG�2�~��k�N�+����5eq��E��B`b4/�u޿G�E�V�2ck�mR�$ӓ������ɻRM��*r�k�O��H7���#��l:i�uj�^����n���n����W��̱�{��z��0x�v
aFh�tڧ�R�ђ�$E�d9�����%��V�N<�@3��qk4��d�Y1��E�oӗ�U�Yݨ��|JXN���G��òVz��a��#;M����5~��v���U�;[P=����� ���%Jf��o0~���?�	\��Q�c��zہ~I�����g.6�������YK��3M\{GSV��aD
6����E�ll�ly�����H@	���#<�r���.�VB��a@-N�O�wU����h~�ŗ������9�
Pz와aay�e�{L�y��1�,�d�Dˇ'}���j0-k�H��l*��j<����(,��L���N���5��uSf6Ǥ��B�$ׇxn	�h�����P�s\0p�#����w�Ia\
�J�I@��zi³�	��4j~6yKc�޹(��X�Vi���!����,,f�i�f�z���������F���)S��oKx� Ńe��: ��](%[]TOֳ�mMzt�m�.�&/��?�.��)� ��^��ѥ�\��r �1Zs9�5I��ދ� L�БjE-�H�D�Gi��L՜�=�����G1�T-,�fN�s/�fg3��?�>����g���!/�A���J=�c�qy@�"jMp�f����Kk�H�R�)m˭��,mp��B���0���RʒCO�%k�A	R?�69��yb!vTÛt�T���Pq����86�C�~����/�Ԟ���I�����ޑ��(y�j{�}�6�b�@W����D=�V��h�cve�)4��`N<��I)��35w�({C�J�|	��ڭA�r��9C�����7�p��e�����WBKu�^��U���{c,�'�m�7V��`�^Ѐ܍$�zw��ڈL��9)�@��U�=���ͩ]`��
��W��ѐ�hI�V7[�2wk�e�#BW������#LP�x�4y5�ZE��y�].~00q�X
�d�'�¢�S%�HtX9�"�p4!a*���i?^�$];�̮���!�Tg�գ�f�4�y�9j�,, �������\1"|����92��P�.UZ&Q�bh��={S��|
U��F��������[�yS�GE�@6Y��8��zk[h���I�Ţ�۫�j����x�m.rԭ��n�톖KE(q�ڹs�[��ȭ^��*��&O�1h�H�eR4�N��8򏰝��^�"�U()�W����Ԝ��Ť� �x{�;�k���] �s7�2�v��5@J+/q���qȂ>0�D��ն@�ms��`˞�TF\M:�-�M�A�ǐ�v��Y�5@!�8�$�o�(c5~�(�U�$M{�P[�i�����q�s��1�����Ů�.9�A����xDV��|�Vp�i䵺߳@v��q	�]�-�ޭ����/̰߰�m2���� d?J��>-� }��iX)i:���c+A��_�p�%3�]���0*���Է��:#c�����MEr܇ �p��	8V[�e�U`�
s����ס1��{C�g�E�r-d{7OI�������{�����/�Q��3!s	��J��T�h"��h����lA��R�����i�r~^5{�0����5����/�m���2Ŷ���ܖ�h�І�kR�i��T*�L��y'�Ly<���*hOME_=U=�;�8��^e��n��o�K�*@�$�lV�0�^
��;��<�?���nk����Eh[����FA�8T@�!Dw���U��e��ߘ��i#�h���
Hi#��E��
�����~�.'-mJ�《ͪ�e�������� ÈY���݋�]� 2��xh��p[��p����Ԩ�&qt+�Uu`SrI+�(^O�Q�<�g�֪}s�`R������+�k��:H��-s��Rl���lcD���(�<����NJ��CſZ���+S���<,�L<�Eҹwk��̶��Z=�*��:��R�f��U�C�Q�,4Z>�&F&^^lC�o&	^�u�j,�|�a\z7�K�<�y|>��@Q�Iu	Ӎ��T$��9I)ᚫ|HY
�I�}�����p��( �䓀v�����B�IRW4���� 2����U�S+�lu�ec���vw���T�^�N�=�â	�p&a�:X���=(�	g�!���Jj��]�i�H舶�B�1�J s�xm=��k��Q�3w��&�9t�I{)p�d��e���P�F�_ѹv��V�`����.h9]I}�B��9b��]w�;� �-�o�Ɖ]�����,�#���Ox& 0��,�Z6VM�?��S�F^n�4*D��Z���P�����^�x���ݙm�o �u�⳸2{Zm:՗�6�+�8���>V�Zl\W��@E���N��ќ&�M1X�E�pU%ԀcG����fA�Fo���'���fȷ0�_�(�BVf̍i���MF��t����ˑ���<�Nnq���0���E�N��y����/;�^Gˢݰł �}R�Jj�LD�`�e�"=C����=�}�B[Yy�%���m!1�NQ��P��fs"[�G��ª-x:d.���{���1�dI�X5*䗱W:�
�|3��0��6�mọ	1�@D$ǰ[^N�L����i�ԁ��'��ج���N���#$yM_e!�ܲ!�C�[�^�q$�w��˄��C�#o�yvVX��crr��H�%�}�P��b2���R� �}p���o����; �u8�X��E�*��q��ЁZJ������F� �G�{�:������*�G�Ƣ�9?,y���lW
HRx��d`�T�m�rN%I\&|v�v>�)����M�A��5�i�cwK.�E�m�&�ة��_�xy�)�����]��\q�֮�wz�kA�J��`����Fzy�Z�Z~!G~4�ş���(|6�穮���F�@�ب�в�!J�f�ٷ�*`�B?��|�e�����Q}�M�9M�fd$ �EP�E�7)S3To��-�����2�y�p��M�8�$$Q�S>�r��#� ��Z�͘cڢ�]�R�/����zI�M92q���P�F�CȨ�.��7D�4�!�`����h���e��i+��g�!�@a��S���q�����31��`�Y�������rB��S6�X��פ��(�e��KaJ�%�4Y6��!F�0gG���p�|��?I�<HN�E�gN�b��ϣH�U�__$_ ��C��C�?Y0��NX�fl�Q���6���H�ͦ|'�n�M?,�}7�n�ai�D��ɘ�y@ZU�U�9B�Qj,y�b���]n�#S2�ƖЀ�*��5JE�~���4#6xn��/V?�r�wQ�HMG>b��������|49d��'J_�$�RV��Ϯ_�(�7�.��w�5U׻z�S?��!iG�OR�E����OE�u�ɜ�qp!��S�dK�Q˞�� š'�2$��Z&}�+�1����7t�zލ��
G%tE� ��6�䋆p<��'�a׽
h��}S��t�F-\�!�3��Hg �8�BɷS'�>�\�c�W�(��4�^��G���n.&����L݆�B7�bgrM�W��zj��=C��ރ�v�$�����a�B����y��Z �5I����| :f,7��5"�.3�rjK�%���f�$�����W�cu���� ��H�ߚ��E�Ҡ#�i�ЁEau���
À;ɨ��{ŝ9DV�mU��NITl�r��H ����A�ϢZ�7g3잫#����խ��t����G4�I�@ס;�L����.�"��C$�%��"�� 2�wܷ� f��r��<9����An�vOߐP$w�`�r��{�]�3��v���n^r�����0��+�Q��C��u�t��0�$�e``;�L���hy�"Gf _�M�����U*�J���OS��%4���V~�9!�C�fз�g�+�y6P�[6(F��2u\x��y��P����� ��W.Z���~���~w�)�����@�%A�3�BX�߲�E�[Xl��M/�x��v��v��&��&-����;3V�)GIE��ft�uK"���ƹ�㑫E�����^N��X�11�ZB��!�=ȡ��4�h���G2n8��\6�u�-llDq\���X2x�Z����6��MRN`�+�<�M������j�ֈ�cY�c^��tv��{G��>�u�3���8��#j����1��I�![q���O����}��,��}�0P��р�?n6�	*��y�&Xw����S�{��Jё�g�pUO�I�A���61�]�DWhBь9��=���<�;�Qj@1���:���p,��(�9�&���\��=��R�N��8,J:rl��$���b|2��(��K]w?�t�y2�ɦ� �j_LV]�q�ռ����,�5�ŁQ���Qr�Tg'7m��C�T@uu�Gͫ�D��D��|i�ETz�o�����~��\�j�wcY�C�#�E�x�:�u�|X���^��:���A�@�0�� {l<�4��
WC~� ~"������]��"�)WM���7�Eۍ�K,�����7H�'oy�E`d�QW#}o��.�*po� e:T��se�9i�u��%F$ ���	�l\?�o�>,�"�h�����,4��Ⱦ����b���^�v�X�X	�W���J� �5;��&�U�@;Y?n��X��OU��
����/a�����ɑ�TQ�Х�aG"��,����X�!�6��m�b˴x0_��M�jy8w���e=��]G�����\���|	�2�2�_�&u��}�(T�lE���=�[�0��T���+�?���iG�t_vF�'�Jm�-`�|�4M�/���z����_�YUt�L*gf�_9�9���˧�)�$�'���u�h�c�Q1���l^�~ǩ��܁���^��-���9����tg��=�ʱ��}�4z�*��&\[�t���֨)�� �l&��B�݁b$��ހ �1|1z�4)Aݬ���ܥ�-�!f����E����,Z,̠�R2AuZ����#��s$O��e�xF{7�ZJW���:�_�6�s�t)�#Ƣ���2L����*�?��e�>�˂�ō5~��f���m�ݼ��~ir|&!����7@v������Za��x��R�Om��mK�E��N�e(5E9�&	UN�Fʝ���U�Eq�<��.���4w�EY榸�w�'�X�%ae��k��-	p�p:��ʵb#��kT�b�ח���/o�{�����Y݄n�wnt��مG`Õ�&;�_��SJ/����^v\�5��z�d�����_��F9�ؚ5ù�0����>qtߍ�Q:�.��n{�L�jg�H�A1CEv�;L�ê�s��M�h�`��[�rm�D]uٲen�PP_kgW[��)A��h���4�{VLt�lM��/��%c�2�z�c�.i�gz������d�j(�=������l�u�� �:�'9\��㶯�����P%�����D������H4c�a�
U��ۦ� F����P�-��*,�Eo �9��ed��}��ił�BRv/D�U�8�������j:�}�; ��u�"�E�r I\m�)��8q�oݷ��(si���i�7V�<X;D���"2���W��;�&H�Hd��sc��mx[�;Qy��>�m�ARGg��`���pb���<E����t�����j_�8׫��dtG< ����c���9�ro��F��e��s��`7��ҟpƂw�==��@�w�7]�a�����r*MI1~��� ��6��?K��~Z��R�H�؝yy�31�km��1�R��Hv^y�~�,f�L⧲5�tV53���9�:��8޵kN���{�����ѭ1*�:��)a�<�r�i�Zy�%��\����C�jrI7�u��{=eqr8(��U�����j���k���(GK௣SR8 {�����E9:2Tˏ�`��\Dk�Ӣ,����T<�c�����n�a�JA!I�S~Ǳ ���9�����o0�{�����r���we������0�?�;h2	�)X��E*��j��rx��eh��T�6�as

�H"ld�^����ф�j�<�퐞�n�&��m3O�9�{DkNE���ۆ��u�'i/&�|�#��~��
�HfF�P�|ֺX��/�X��N�_B����W��)�F̬�cQ�߄�r���[����[�#J���0�9�F�m����gY�Z� 8��5�엳�<�f������O ��ǕOā�~vh',�a��ىhQ��=3�=h��9Jb�$���{�vH�01�-.���M�&;�7�gOu�����_e��<��(G&j�n8Q�d4����G�\�5j�A!���f4x(g����R��;Q�C�>T��S�$pXU{Ȩ)T��XP����p�7�ߊ��p� (����?�yK���U^�� �?�! ��ű�"�pq;zs_+�+���W��z��0�0�Q�l�(qUV��� �H�>M��,����$��x��`����~}پ�Iv�醵�����f���[0,y�'�1�B>W�m��b�������Gx�B�S-��w��3#�����P���1ˠa��a<�O������KX�kt�Cq�05�I�3Ի�]���P�>1�9��"�%�:��XN� ��3��	X��A�@8L������z�6+R0)5Q+�w�j���A'TOl�!YU�j�ଋ遙���r��p�&t}҄��X��uM	l�5�!̠:R��3�ڽ�������$��]����<4���R��I��^�H��T�����a~;����d��1X�hl ����jH����@6���K]�P��x�����J�����>��40���1'QŽvoD�z/�x|��ɕk�ԱE�&�[bD�#ڂ�g|nG`�����W�3Е��ƭ���D#�Ψ���:�sU���s���y�'������m{�2&�(���9���VQ��;� �ΓB�IC�f�����$T���p=�R��l�Z�IL��*��w84�U��'ZQU� \���Z-vi��4R�T� �>�(l%�����o��W8���v���ܴ!���C>�!g6qđ���e9�M�^��$����� K��E�{��$�ڥ3�ܵG�RrbE�[��Mfꐃ�WbKW�(hο�}����F[d��Z��.w��y���D��i��S�u��\N��A�ڗ��b��?|%tb���^9�@c��_*�����]��P}�O�#�-s�~e-�@��J,!MN|[��*����O/Xt�Nݮ�~����[le��I?��4K;�����-����� �~�{�Xӑ�Zt;�A6�^'�,)U�#�&B�[}ݺ�jl��D�~�A�RbnZU��8�CJ��P�λ�iO�С;>�4]�*tƘ�}5b�f��Sn����h�uZ�<���S��:S�� �*Z2'���i�X�W\�Т��T��ܽ����l=��e��ss���"[�zK���`�%�`�w�Ř#�b7�w�o,�K�h����W~?l�t�qD�	�c���/@Y���l�m��ͧ�܆�?5�	���Q��8��C7Q-�eE ��f��޶(|Ut�ح/qDH�*����`r�"�AƲ��U�T��rl�ʈ���!��9�C4{��r5�����X
�p
ɚ��q�����m��ڢA���	�! �o�˯��-
�$��V�&�|�9o���,s�]n��f���4k�pӅ���	���F�v�Ҳ)}� �Yë	����s��dE�*K��U��� y�&��$�㯗=:��M�)�D1��%���Z��K��F�L��+�ɸh�ABJ�pԉM������zysR���PU�B���bN��dc�j���*Nƛ'��� QQ�"S>�l!�u�Y`j��A9Ǔ�����ol��cܡ`~`�-�Jj`�_L5PR�`�M��4�:��ϸ�FI:���e�������h�A��p���қJ���I��ڭp�2�l7�=A� �Fe>�ˇ �B�7�?�"�1�y��edwD�-�({W��R^9V�C0wͯԫ�Fw�jT�8DgI�-ծ�����q��W�6aY���1A���^�C��vH�2v�t���A/p��OO�]�U5CZi��>oeA�Ϡ��l�O���? ���,����S��z�zع^	�R>2��M���A<�4�A�91x��>�UD�� �����|��\����.�
G��.)�~�p��&\�D���,����`�R9�C�L��8/{8�o��U�j�B^��Z��SҾ�U�Y_�	�	�(��.��;l�]2�n����+d]	93(�E,�/[#7�?\�eA��V��PK��W�Q�"�[���(K�n9�^fď}�b����q�� �G/r6�Y|IE~��zvF�����_b���6&a��x���Im0�֪��]�+cڏ�z=��Uf�!7�r�������'�F	7�@�DIƯ@�H�­�7�B��{f��8?J������^�]��`��!�[��q��f��雯�������H�s�Qp�� &ߖ�D��Z0G�yc�@6�=����?���X��d-��T��[�Idm�ѦA����ڍ�Z��Q^d}1�o�gM�jn�&-��b�D��68��%'-s]%���T�.�-����V�гb	⊊ �lp�>6t>U�i% =��@,�X�B��=$&�Y��ɀ�4�]/=��=�,q��}��/I%ܥ��sr���}�42�n55~��ΰ�E=٥,_��M[�a:`��Z�ܯ��`�������PRl"�ig�E�:��y�/�����M��H�V�e j��H!ߎ���*������Q�a��@�6LY�d�2��d�/�F.�cÄ�
�S5��_S�,�����e����B}�J�߶�j
��q�?�Nf�<��hw���I&yy�u�x��H��w��N�{���v�ͯ���k߭'�W�mP��Lp?���d0�d�M��Mˏ�|E�
e��e�������JP0'�W*���|�����R������uW�A7�(�xt̤���}���́w�-����������I�Of���J�ս���Rĵ�+�E�5����)����l��ѕ9l睼':�?�Bd���M��Ӭ@�/S<��7�����F�3���]�^�+̗�G4���}�����R�=��y`2��dQ�����39�΃?S'�g��`,��·W�b�HzdgFP�k����=�b<H *�~�<q��.>�_"�Йr�E�Ȇ�� ����Y	c�z��'r ^I-�O���SMÑ���vx"�J�p���BcI5OT�%�	�,��30\��eLA�x{7ߦ];N|�/�C�'D`2�t�o�Cmʼ��b�m��]���X,��]�c���䱟�D�� V�59|\]��[Z��N�TX��1]=�j�ǵF!�7����KQuzM�n`̆�!:��3����{+)�Xpf"YF���;�����B(����@���^�4�H�i��b��Farcd%}�@%k� �����e��4��2��^F"?��^
0:�m�%���_��� S�Ⱥf�0�m��<�1�:"�]�h�({��v8?E�pH�\*Ơz�*cp�٭ǣ���vN�#&�R��	�=ڍ���!Sy9�����=7�
��Ff��`U>Q+�K]?uց�T�l!s�����+��^>˟vn�����y�������f̹Ne�,e�R���-(Y�[?a;����DQ�3�z:�={�oW?ף*ك�t�7s�:�~����*�4
1#i��=��nnΓ��6��8��s�m�׆�@�nԄ���Fwt}aYQ0!��K)�d���l1�l2�������ʐZ$��;8�{#wf���lٔ*I9�>�M��?�?K'��7��YX0e�`FY�b����N�/6�2�!�DjI�Gn��ikP���=\F�r�f#��]-f�@r��ŉ���~/��Tϐ�t�jT*����qUU��I4�2� �j�p�E$�`�b�����$����`�V&ٌ�A2��>��eAw�d�ۄ���ֳ��{�_�n���y�Ue����S�~��#��2LD���(,�tW���A���ܿJ������������ȴ��
�%ZA�3����w�K����P��S&��@A;`�ǒߏ���[�ĥC'�,]����]<�8�+6p"�Ej(g�Wp"��C��m��@q������&r�2���	�Ϩ�� �o�ua8����ǖD��ٜ%�(����2`�b�Y��U�U��Z�{��W\l~o���ȞG�]�8���0dܱ`�m��_d�O��:Y�����H���xyytfG�:�����3]���v�W�E8��ݥ����Yt�خv��S�<O�KD����[bҷ�U����};�2o�7�`���1����k�;���	Y*�4[I�[Mp浮8�?�h|~��d-c3բ~�Bqo�Os%���ϸէ�n��ߢ�pK��B���5tx��+�{
��]�<$��\�+"t��/E���UV���2��:�,���{Y*:�\끇����j���n��yMt.�J�"������)]�L��>U�n�ϵ�'K�K����z�gG����|'���f�D6ë.#j.�q��pE���|�R����+:�h��$ď�-3���BpC�n_��(���~��;n��[K���\��.�
����RUjY���/rn���_�HV��`�,�J�:�j���!ք�v�J�}�(�A�z���Y��:�N�:�S#��z�,�a��n���o�%��}� �NE���(��'�Sin� �.��p���,�M���m�SN�n��������Sc�Rgf�{zb�;9�&���o��BόV�'0�
�=-�#�����>�9{��U�L�� m������?g��bnA�����2 ���&(����I>���g��B�82��5��n�P,D��C��+�;���ģ�*�r��:)�n���9`��v�!]�w�@�-�>��9fک�O�D��(ϵ���ڙwW��f����5hg��e)Z�'�X/ ��i*��~�Ĝ����3��u�F9��ro[��-� Z�+"��f�"Fsk,��'��v�u���؋lb
!�e�y�}c��$P�k�0�����x�5@_�֨�U��N��4�:��J����8u��i����}�~Y����3��~���	x�qO$ TB��c,]�V���7b�p	ġ]�h�u=�t6)HP�"b�*#�ډk��=�KM���5h��o���~s���0��)*����'/�p��e�8�}��<�zc�bM�F���e֝X��g���e��hP�}~�������*�~�B�jm�����V`Bo0�=��GU�O0�VK�>���Q �޻V�`LS�{�h����E�Xcj�25E=#C���@`©'n`B<݂��F�.A���t��y
������l�͈����L�4�O&(��zє IԒ6T������Q�-����kyz�, %��;�9!(ɤv��k�z�`G�T�i'��U��G�[�i�Ғ��F�WT��^����4��=��)o��x�5ډU�i3���G,�EY����HN�������2��۞d��vH*i��hf��Rk��P���OY�Sk��**'�vY�n�H�_r ;�+Lcc~(�e��*�[�� w�(gMr�?�<��a��]�/!�w���,E%l?�1��/V6r'�i�~.K��y7�M����f�
�7��ӡ2w2)���42j��:l��[s<vM{j�om�uOM`��W�\�E��i�@.ow��hp���ݦ&t�\����-7�q����H���ũ����� *��޹�6�X:~�ө�S���B9$�Y���D���P���Ո'�ǯ��~Km�L�ڵJ������>ܟ`�Q���!��.�uRQ��.�����Ž3����s-�!o]+�� w �e'�H�7�V+�Q��ݚ]�sA;
��m*�RG%7�>��`�%Φ)Yg�?v���A/�;iG�DH$՜��m�q��S!��Ya� �xVgHH�[��E�饏����B0Q�-�RL&C��B*�ƫW>�Χ��o(>Ђ�f��	7V��c�%��RMt(��>HVj�[��X�*sK��k�q'ӠM+Y�C7�=�41:P��g�8s(j��F��+v�A�\8;���8�?�qG�2�%n�t:ך��E�!����RI��4�yS���ׄ��Fv���;+-�"N�VJ�����L����8 2eil��L�>��dX	�+��W�}6:� {�:^��@z�����AO���ƀ֦�3���1��YJ��8�F�.n֟�O�hn��w�}�a��~��kK�����������?�W�������F��f����Y���|�/�9���Q4�`���@am%J�U�t��C�A�?J�ND�(\+Q�,N|���O�#�ǺrM���I�C<�f�6H%�<��b��(9rQ��o�4�d<��s�����t��^Cw2L���Ӫ�?lP�(�/�����ݶ��9����T������o���Gy��J^҆mC	�O
Fgl�s��3�g>Cٵ�Ug?�a��]��`��mSm���N�ֆy~�f�`�ަ~���4)Y����M��� �ǡFMI ��f)�R�T���K@�,�W����^R�c��Z����zp.��g�"�*n��d�#�qp����Q^���_��G�N/	9B�YS�b���V��QX2;_��ڀ}�\�'�A����vL�ˉz����&,�6�_�ge6�!os�!����r����[���WqE��y1��	` b5�ŝC��:�33�c��A�>�j�����eC�a�3��s�f���z�s�Za<SD��؆w̚N�j��^�a9��g�A׋e�݊�Т�N�P?� ��Q�J.\#�x�'ui"T���\��7Kxʣ�NE|G��lN!Փd��t����e��_���J� ƥ��"�g� ���"�uf�<�ki.Ȯ{���n� �F�=��ᝄ%�.�a����������j�,��hɴ��G^��~R���2��0���v؉V��aa��Ɍ�X�P$�*ǟ\\1��о�51�����0�c0�ţ}ZE���-�_���lQ�F\ �����,K�~�R0UzHVk��~tP�3����fץv8���4�fP�}͖3�}���bЮ}��w�M���72���m���T�a���0�	0f�w�Usf�[��c���&沒��5��s(��̠�dq�犙g�.a��Vh��7�ж�8��vS�\7�\#���w꿎A�=���\)�Y5-^A�`���vՋ_���u�p��J�3��VS�����9��B%�'^]t]��z�-_�X�^�
ψQ��D���3%8	��?"Ǐ�f0G�h{�8�- �����	��7�j��q����=_gD\�0F�Q�C5��d���J\ <��3d郢O{*�4�*5�3��[�2���ǀ�C�E�T��A�}g��qSY�$�VW��xj�]���DAL􁵃�Mg�}�此�:M�s������+
�H,P1}	���砫�uN�M���1	k�RJ!�m�м�r�D��X:���^t�Е�	0Y�e_7a��l��e1�juݺ"�=��u�!�T@����fTtO���fpsp��|�n�#�@���`��K߰8�(�?�Y��ښ����,U�v)�N�W�a� -OJI�{ܬl&����TB2��_�:���ܺ������cd�RS��W�cZ��`��8S�C�!="�dh��
W:ݦ�.{��c�1�N5�2�<&�(�k$�A����'�ƪ��������U���A�L���)���_4(��y��j��Z7+(2��$��M�nP�~8k��'��b���8-=��*�!Y��˟��d<0!�ǭRj(7��gh��Ʊ�ᣌ_�+����۝����nXx�+���Y�&�����ڻ�����b�kt�X�-���h��'�$�U�W�!_N��m��2�&�b���<1�+v�]�;�#�΂� �EMMzBL���[S�Y�?�(����UF,`�}�D^�8��0�Aڥ(G@^����!z� nBa9x��d���G?@��Z����� #����q��&��G- VvN�	gb��JBK�	�l�=Q�,�M&t�-t�9«�M�������FN��^l�� (7�z����O(��[�h���cU2�X��.�h���@:����Gz�S-�d��Qg���r�4�W�?@������m=b��."�2�Y���I0ab�I�����c�
�4Sn�l�5��4��ᾝP�[~����s�Y�Rh�$\RC��Sz������u�l~C�؎�h$0-��^F�h�*Cx�����Bnq�/���ap&��0���y��ֹ9��x����K)i�;;{<��	0̫�w�&˼,f�{����
��i��.=����u���?�	uA=�,�3v,�k$���9��5|Bvhq,�J)�/#���V*9��M����T�\és M������_1���o��K9�Yɜ�wa�*B��1��#���ܚ1�,��:����E���2�P��LRب �یXg�&b��He�z`��V#��i��I�y�7�NF���)�v��o�
�Țg��Ęr�^>9[b�����);�U�v�[2�R�'�o3�>O�-z�U�����T~/vf�U�Yh(����q�e�t��3٦��#�v���=k~7Y-ie�E�����}�G�e��g���/�%n��&,�j-C<�C���p*�lb!��JS7��`RLIP����]�B����{84�喏�� �O�炱T��7�O;�@�P7�źCjNC�&.��M�[)U;��q��yE��z�oa{6�	�bCuMPN~8Ϧ�U�/D��7�c)��ũ���g���S���O�ҘՇq;}�o*����d ��\j�M�F]�Xr������~��p5릫n�ovp
/p���bb���@�F��ʋ��S�T�F~��K��s��>K�@ߠ	���.h'$�����\W���;��~��%nT=�*Rv?1:oOI�J������v�T�%<��&����cUX��$��f)��t����jW8��~IrԆ=lC���f�C����R�)&hz*�Z�����B%w�a���r(R=����2��5�I+�ks���R%�a+IRfM�G�B����5�$�	?�n��ϕ�}�T�^Z��eYS7$[��}�@'��Y<�@�ӽ�gS��}���<\�ɬ�Ꙅ�Ѻ23;��\BP�*ʨn���� <.�"���-��A����jw1��3+���<���m-��B�/b2��W5��]�P>v#��uHfB!A����d��, �h������`�͆��@Ai
���|ɪ߁$�p�6���������E��E��p�C���E�����>g+�K�8��ԫp�8T��+�����.�+�F�Sm����1�������.�&F.�Vhs��`�0�Pq�U��N�~��U�Y
<���O����V���J�#qAZ))�8}qw�.suV��)�_�X�.t7c�(W�*�M�t�h���؈����$�����Cv�"{�7��\��Q��) ν��ݕf�2�eY��Ern�������+`;�J�&�NM3�Wl��9bJ�|������[y�!�B��	��>�M'o�)f�/r2;�]+�sm?��/yO9/���U]�M�V7����-��M>�ch���E��J)~��Y:�?�-u��d���w@���ƃ�g�R��@�V�5����P;v/�e�]!�B�E8>j&���D f��e��r���RL�������B��z�ɢ�E�G��s
��������h�z���	��$��t� ��mqU����\�㫖8�vG]�4
�J�W��
��u*>�Jyt $�����$��o�y�Q~x��(���5e�+�y��Z5 �2��|�D���p�)�-��_6�=-`++�6?<f���C K��H�oDj�4��n���!ވ��QT�yw���Q��d�`S��z�g��S����&K��ƫ�i�A��R��:����-e�^"�eڊ&��pN�G��+>�%���NH���k퀠��"�E�"����w���Gd%�]��YS�(0تr�[�s���)�ա�**�K	��FZNP�Myɇ0��9��@���x����^�-��E��{ ��෕��B�-��وhݳ��o�6������X�7�J�%m���	��_GJab|S�>!;�{NL��|(1B}_z���Q/�L>Z7�U���I[/���l��<��l�e��E�uѯr��r�#�[����()U��vY�d�����o=��p��-���y,������f�2 �����	!^zttDF��*�F�ײL�V����&/����wF�`����/�k�p��/����r�������-G�!'�=O&�3�M;�a�Fύ���'&A��p�(���)r���h�Qv��il�A�-��}���Ο�����FЉ?�̆���	���禜�ˏ#ͷ��y��D�!�٠V=�\��Ɣ2��vR����a����k>		�)M
� 6��U��e�ï�1l��'S��|�?C,��հ0��Nd�)Y��)5�g��`���o�k�7pX�]������TТ]쟞��y!Ô[v��Ww�z�����]���+٢�ѧ�+R�)lu��N޴���֮�s,2C�$-�'�8qD"\וc
_�h>�W�-b#Y�1��7HC��߬;ݝ�����|�F���+,��*�­��xno�&�|�4,/�x��Su4G5s~�wV�'�)�ii��Q*��S-)@�Qc#2)V�k��׸���ٸf��K?nQ5���!��N�°Pp|���7j�I�glaZ�������f�Fd�}V%(�gDM�3?@<��������/�s��[�R�'&ڄ4��g�i��~N�h~�b_�G�>��`�]�� �G.3�|f�ga|f�}��YȊ��D0��q&��/+�F�cG�b�j�ğA�̷�(��-3�>�q�ɀ�c�*M��L��pe &,�T�R��lW���6
ϵQ���Cr|��e�+���T\����u��%L�@?ā�/��TtΓ�M���*�Ż��Cqı�+���A=�`*�[��o��� ;Pd2��S��Q��!�&���\��y��]�9FD&j'�)u,5��rL�BP��])҂!_�+��amK�)ĹO��xEu���Ȭ��桨R�8���a��{�9� �<���f�ȽVig3�U08Iw�so�t��s��Ӫ�$IM2YdQ�A�N���Y�bOH�d@�x���D���q��H4k�Z4��V��x�̪�WEV��E:>��6�Fǆo}os�)5M����I�^�6��9��6:����`D�6{|:���S���E��y(gN�?u叚�ѥ	�Fx�Qa��xJ24H���sX!�NM'4P�B�~���x𯼌���g-�~V����Ҷ�d4Q3�Y�8��c%Jmk����Oa*Ϣ"�����$'X�����z��3� Lf%�0�6��O�D��g^�FȒ�l����?��W���<�œ=`��߁�g��k�[�8�.���O8�����0�֟�إ%?-��G�:26�8g��`	zW�-FB��c�����}��ĺk���
��_d7��Yvͥ�y�g޳���K)):6@�yl}/��P{��A�}����	��حu�
ط����3^U���K�m���[Ҭܵ��.�����5V'S��UY]ag(�SC��*b��_E0�GZ�����d�9&�#�/8�( TR����;����_x�RD��B��d�2f�Dԥu��������/�K4��V��r򰵚7��yyW$ˉ��u���ゆ�w4c��^��d�&n�7�$
y�S�]{��lY��[�DI,��`�1BI�н�d�[c�;L!nz�A{Q�:��g2�������A22z�7�kʹ��N�%�uMR�����;љJ�B��pas�����sw/P=����U��
m�rh�ꭹ�E����K���o&�Xd1^����?q��a��[;��^ ���Sg�fB$lsbS2Ū���(�^�V�Z@û�|<���Ղ%��:��h�S6'��s�·�:�b)y�O�方�nt�j$+"�������٘�S�28[.��5������`��~���2奪}��C��;�KzM��l>�m�I�ݰP�S��Y��FV�o�i~$�ߔ��,�K����5�X�1/Z^���䒕Q��,�<\�9*�����٢i:�R �����^��~����DM����o���"@�z=��I^��[ T��Ħ��T�Nm �i@v���C�!��Gf�V�e���%�e-{�D��}�@A~���,�d�/�y�0�K�{�<[L�4�H��Eg�����E�1<И��>=q���=��߿"_i+u������}��0z�}�L�ReS�T�PD�s��&q��������W�%���M-��J�?(��,�Ae���x]>2y��ռgX��-	:�J�t�@��*���r��`G!��%�)�@�ksL���Ww��3�j�����qݎ욪�r��� �����ID�7�&#���e.��e����tU|ˬ��(��@�*�|�9��#����q?���RL����%���t��i��d.���-޴��/�����*�D>֔��Z�H�9f��_��v8"����"&�ڧ'���Y�thw*�D,��l��`&�ޘ��%��z]��Oۻ�֘���~�I4m�וP#�DyS.�/$����&���46i��>f��ݙ}�?C}�M��<�+�m]m�Q��%R=����s�L��ESxU�_ ���ޒv0ot�\��~���=J��&6G�� ��B�ޏW-���Ůs�)��0��B�W�``��`K�*��6r:����^d~d[��*h+Azi0p��/�|ό��S
]�(q�)�۲[��5����'~��r�ko����i�{qpY�|�yQ\����ڡ��a£�6fݾ�?�.�5�*�ʴ�q�ql<���{1�`3Ǒ�
'�G�4Fq���^�W�� �t�!y�q�5=�K8v��^�-���0g�_P�O��T�Zc��l�W%4�	��H&3������Q�N���>dΝ��UP�����wk���r�y�8c�霐PA��s��A�cu�B�6b�g�o�,@mf���,,`xQ�J�mj墮�j
����Fܗ>��^ش��XV̽�1�#�j>L�ދ�!��K�fa$�f�	�͹��;͊�ͤ��?%,�.[i����]����-��)lM;"��
v?x��h�wIvk���!<{��
<��=[<f�h1���~���7��e��|2̡*���yU?���ER���z)?Atp N��W�!����8�� [xj�����'Gq̙
�H`��JDM��W��Dk. C^?���R�60S}s�4���I�����������h(�m���Έ�v5�V8p�f�(c�P�8W*������uBu�6�t���Zf�@��b8�<������h9�w�v�ku�>V�MI>�&���5R/4#����u�G8�
���[��A_F;�H���5,��U�>�ٍ4�z��JH���M� 3�b�����f{���z�z�����vn�R����cK��!'���y������Y���<CA���7#�R������Y��be��.� �.Ŀ���C*L��/z�D����+�b�.K���Ԗ���9�h��"�eG63>��?������E�ǊC�7����f�N��÷�ci�\Fw�5��td)Z��M-j~a��o $+G�V!���˞[h�c~��Q�NÔ�;U�0�� =�_5��;�K!vW?K9p����'��)�ܾ�%
��כ���{p��欶��|� B�+l��A��M?���>4�	`��:��сC���h��f�;pH�xK�V�?#:��F�p�ɕ:۶���J�78�-�*�5�1��Q�D[O�*�*������O�5��N�Tb
 �j������慄��p�b{i����l��^LG���j3��y��V����Ux���|7�O�M�偌{�f@ŝ���2}Ykc^iE�0'5B� yE7؉۪��s�4������@�YB���O~b����nj�w�	WW�	�7|��Fao��S�H�M�v�Ȟ�bά|PQdY�|�WS���VG��@
�,�����F��t^��|��4{Z>�1AnvՐA�*��h�O����X��5϶�&���s�Jc(�&\1�GJ��/2�rNT���
S��Tq��0

�W?M����R������,4����/P�(��g695�I�dYdo�i�xqn�����NtZ]N�)�c��%6X:�I��o�Al��x+#	c����S6���|L�,1]���))]we�&Ҝ��nrv�� w²�P YO��if��T�H*��/�d��Oʨ̯�-4�ke��=IJ�y$U��{���%�
/��8W�O�ޮ��? e
���>>��QZ˩h�|[& ��~5��\���H�z������yte�쿑%����-&6�5���<Q]+�^,�{���}I����h�o�e>��W�F�H��3�/T(�����d���Jc��S�O���*+>1}#�;/ bv��?�W�xn곎+�U���)��,gJ �4���.�:xl�����'�/Sby�	�R|}7`���.6[i������m��ҝ�S��0�#bU`K�tjK��ʎH׋�.��~0 ��n[g�0��&���^�ץ&�QI���ގ�!Q�=#b� �{X�j�?�SpvtpZ�4��78��8�q�����h���5  ���G�M-Xs_1=�@���7t��<Ds��/O��PH�T���[8���ߵ�K��trmu�������3q�~?���2qcK0�EI�m3��if`k._%�x������V��x��ۧG�� ��I3{
Ӎ�,Z͌�f��alz6҅���Ǡy�M�4�R2>���D郀�����V��k7��cw@G���^r�ͫ�By@�e���������H�;��E3j��Ƈ�$�f^o�'�G�r�^~|�h�)Bu�igm� TZ��^�u�v ���:)��p�,�8��O�S����R��V`�e�?WR���89���Z�Q:x�@��=tÃ����)�6�/���|��S��Ʉ�ܱ��}��u�o7�³�O��6PUaB<�e�����IX�d��,G�9�~�Wj��:��Br�CT�mN�7�D#?̵�H2���m�YW�B��,@��=���Z<�8������M����y�������������l�#�|��iwV��	d���t� s�l��p��	ő��\�Q	�v=AVw2�4���G���`����ۦmR���PKA�Zj��-� .�������zҒ;?�,)��r�T�wȉI�N:ht﫵�4���T�H�v���Wd��Әf�u�ݩ9��P��^F~����pc��7�����.�8�Qil��E:f@�t�3G,���n��;�V�6˝#f��?����'^�Q�����q��L~\T�7[rF��,$a���7�R�"
��EϹ��/2^WfaE��O2y�I��AF2��
(�,C�-�e퍽ܧ��9�Rf�)�������I�����:
��t��Tg�,~`D�k���lZ������D�ņ|�g���~�6(o�q*pO1����Vǯ~3]��in�����g(���ID�~�Z���@2�n�}K��%�Bݷa���Gk�om��ŧ������Y�]/�Z5/�g��7�����cB0 |�<,�R��H�:'�p@���BGC�,�,l��˼�v��H~�C��]�D����mO��C��V�O�_BP��n�F\TӢf���hK�Y��]��`�0�䬼j)�"]�s�f=�R�	g�S�hd�@�#�E����g�#'&�����ITIF��ڍ�J�A���j��5�α���KWK�vt��a�:*�8�'Y`Z��f�=���7}�(~-r�B�畔�a��=��J�:�P�d$�j����6�3��>J�X$F�m��8��b�t��V �]U<�N,��ea�ޖq���P[K��R&�V:H����hO5���ܷJ�~'���$5e��;�����ݚb��w�"Qb��oʶ�^2������%	�T���{t!:mm��=I;�y��mP��"k �I{%HPUl�(e�����y�o�,;�7,��l`e��.w�t���F�&83q��0�c���4�����
�r���"K�I���4��=�id'�6V��?J
��ŷ�b�	�1������p
0/�����+�p~,QyXn�B�R㣷`!�5W,7�I�GԪ�cJ�JK5���=�cv�&?�֯Ү ���<1�=1?Ee(OT5Fɍ$���#�ȟw��Iݲ NC0�s���s��
b��`�$�a�I.���e}"�����I7�@�j�%����c�YfVr�%m���.F�2�5,������i� �5�$Z���E�u�i%k�7d���,ؒF晵����y�\�V�t̻ص p[#����9;J���xk�P�A����k�?��B��W�� ��I#�u�9���U?��m���c��,�UJ�P�1�*!s7���Fc$X��.1��#F�= #췚n�I�]|���dX-�Qaw�����X������UO/�:�g߮>`��צ�G���V�������	w��{ź�E"y����/Eܬ�adeCY �<�]�{��8�Jv�ԖN"��p('i7�qs(Ra��OBT���d_�tTƾ���6��,O�?�m�-��gӟ���*����nf�C�ߜ<r�e
���� ��]ڷ����M�2L*�a>$[8p�UѲV��AqA����N�B���J�'�:jF�[D{����"ˢ����C��}��"�_�;�t��ը��,�+�؝�������.�,�w�cE|�n=J�r�=?��K]Dv���+>��3�f�6�J��ĤE}��ǏZ���̰U��5�=�R�N��q�^���E�0��|���.�ٵ�1;Sw��	�5�yg�w����\��6�����ʳi}.��e�I�'f�C���1���4���ґ�a_�y�ASy��<����誟ֽy��@�1ϊ�l}��xf3{-��Ű����������&+hN��"��3<f�J�d�&y3�',1�z�_��2,,�!�g��V�����pE~R�]�S%�-Lt��V����\�S�����-�������v7�&6��B+�Wr�0�s$
�}���Y��b��kuy�hL��-{�����J����b��!�!�+��9���O�c�w	��	V>��i���2l5�t�(
N���\��({��8����4��ӝ@R����<FrD8��m)-/�J�Ӏ�Z����+oH�O�e����:q��⭸��ۮK����A��q��Y���f��_����Ǟ�5Rt�^��s.��b�?&����Rn�_�����/J��呍��G��h4oߘU|1f����K�컥�3,����J]�</���	�[�ڮ ���>�ٟs|��B�lO�} ���*��4��}��얹|�Wl4j����ל}�[+��=C�p8C�
�S4�?Iv\�����Ѿ�&sH�&.�T��s�ʘ=�*�޲QS3����P�rDlm%�X3�[�W�ŧ������Y���_X�I�g(�P�aL��m-��>4�0}\���uN�P���%^��~��z�sE���Dm��!���2�l�?��Ԣ�hT6vvF��2�!�Q�TF�? �$"n�Sl���1'�y�(0���,���ފ%J�dZ�4ҿ{�-n�'Z����6zt�����p�q,�9�p1i��ҁR^E���P��Տ;?*��-��1F}�"@���j���y�Ǔ�G��_ ��|�ҽ+��a:�O/B*�u�{�=i��n$�!@��fK^������R���F�����"炐q7u��3`��m8sV��BTh��9+c����&4�������=9A��艝�]���k#�f僱���y�;��y�@il�4�w�vKy
@g�?!�FuV��c���%fz�](�}c^��r�x?k]-��h���M��P�;x�|��V��/sJe]К���p�� pG:�
w�8�ߣ�dlvz�VZ&��=�W�S���;�����.O%���"�l��x����3�]���uzݥu99�@�L@.�Ƃ�C1r�k����._m-aꠡ�.A�-#�Y{b"��gs㪹�{�Ǯ[��T֯�����+qY�����I�!���ܕ��*jg���%�0זZ��S���h��:|"�s�ݙ�ķ��� Ob���su=!ϥ�q�R�78��x�����|�ڔlfV�����e���+S����"��v�.;#�O\MaM��I]���A9��S�w����@��Z�*3�	�3� &�t;W-4W�	��M��G�Z%1Y����J;>i�U1��~���FiE��+^xn\�d�ײ��--�f�%�WFJx!�����x�4Km��
�3/fh��wBњJ�U�B�7r:s����Dȗ:\�<u��ޔ>g��� O}A��M�pe���`vC�$rf"G������3U�U^���{
%\
~���8�q��.6BG+�j��Wo阫���j7�d/KK��&����f+S��WK.��}�ra��|�*_v>V��4L�n����z����"��EoZ�����T��&������r.�(�z���]c�»�ו=^�bV4!�Y�|<���g�1q�;�4��+�`uɓKR3���7������锗��B�����E&ݬu�S��I�ĭ�3!�Ō�=A�1��t,f�dnd6�C��5:}w�������}�~r��%�{���h�7��ڪ���a��P�a6��+��?�G�O
�-Ndyt�޺"L\��D�:!�g;40���@���H��X��{q�`��3�n�u����H�F�]�3� �B��;��� �.c��9��M��c�a��ٮ�%�R ��ۇ��e�,By��\Gv��k�B�d�:=Kf�6j�;)w����nMYV���5�őM�^�}��Xf�淚��&��������B䁟n���Ql>�����|�k$(��h
�PuDk\��H��;��bE`3�8�{A��z����-=��_毶/������[��BC�V��ʨ�1(�کQ�ϏU�~�)�a[�e:<�|M��n�^ 
�b6���*�2>9y���i�X�Yf�#$A 51=� ��2��#)��&�6�+��'��@������_�q�ٙ�!��(�5�U��T���8|�#�&��6�X�u^��1!Or��V�:u���k�Y0��"3�C6�\�7���9d�p��ڒo�a�[&Ѝ��(F�w�n|�h	���oX�㡄*&������C5��xz�@� G2s\^�M�6Dr�VM�J�fW#g�{�t�I��QcQ�dR3�o/�
H,��b�	Њ�u����k�*7�_d��3)'h�H�S,1��[��������nvts���c���AT�h=�^�C��0z_�k�=��>*MB���O1�s�/�kV�it��b�jG.�Q92��~��(�P(NZI ��1�.����Ě@ź%q�����w�3��&�
�Gb��-��g�P�l�p���F]�2�;4�wZ����=S����$�H"��hw�$��W���ςm9K��Y��/�OBRb�|��%�i�ИG��sE���S� F���KǸ�/��I}�?a�4F�C����ߓe�U���z���^\��L�N8�`֋��� P���"�����z*(�&n[C{j����fpN�z��Ø���'e�%��!H_˵�W���� ��n��M��v�%�=�� B��d�Mn�ׯQ���M.��`Uݭ��c�z��;%
�r=�
-�MV��2��^�� (F���鮩�[	1�#5��րB잳�$��ٕ:ÅI�4�g�V;�1u��=,U0���=�F���|��B*X +hn`7��;��q�@�,l�ލ�9wh0���}�����D����U� ��D�! vR��ls��D�K��Ӳ��*t"f�Ƹ*�����V �z�z��n]:!te��8��_$�(-O�z	�CA�1�s�BW0�Q;�e�q@=(G�H���"�W�6G�8��|<���uڬ9I�r\ZP�T�D��	��S�~K�ȴ��;u��P���z(E��zȂ����z-�fjoV#����iU�EV���б��=~]�<���}7���G�v�/8�r�G'��VQ�*+����)8�6�#�����n������b^ɿ�(b��(_x��2��'�������������Ҳ��XI�j?�<�������7B׋�'�;E6`K4��L������{4bx����Y�5��V��m��4"�������1�x<A���6����2��}�����}2OA͖z�ˡ���	$D����T�s9�y��B��(JNS�K�ZJ� ��+"�eŕzZ�	�r��d�F��8�#c�����I��&eL� ��j�SQ�t���{6x�o�����}n�58+���X���<)5�/7jL��З�~p��B���-<��3�/g��
mW@��|9W`[�(����v�'VM�QR۟���3}��8���l�o�n����:�qF���M�ip��� �&�,�a�}�5JN���;L�i4���g�(a�1�#���gZ�ԫ}$��zjI��-uɇ���Z���,R�L��h��J� �	f�OZc9ۈ�t��
[;:Yν�ռ
�12��7����gQWP|���v!��AF㧮Q���i�J�ߌze����:yI
��_X������܊d�ݦy:�w��~Jx=��F.�Ŋ��8�fR�/��
���G]�mgH���WC��?�P���|���gz`�_ǚX
;+|����<}ef9%8'g��r��|�>��^���E4!%>!?�)�qw
Z�Kr���iz
��ݴ	{�PQk�ͯ�*f� �Z�&�Qd܏@�G�eU�֦.N��$�0���_H��J��T9�1.p�\+6dў�o�T�ȣ#
� �?���~�1_�(���E!��Է����j������on��4�M�������ƍ�K��#.�n�~y�.�{�N?�|�T؈ I�>��׆��yꂰ���C�U���۫�ua�!4U��I@\w2m�\��?�;�8�+z{VjVX��I���������ol2������R�#$Vp�琟�s�Ɖ�}Y�G���i?�k=�� f�/�`f��N�����v�����G��K�oh�xbO�&R�i� w�ЉV��O����e�����h���ˢ�e�A�cF�
6�2�F��	k�����}�kHT�6sRmТ�0^�dZ+���|f,�S����E�$�1	���'d[yɋ��1g��\��k�� Մ���SV]�"�q�pMƥ�L���?�4����e�CKXhi����~�"-ڹ����53�2/���s��̲��|Y�n�s�4�u@j~5K {H�6y�E�z��b9��)���m9r��$�^�H^tR�k@�1��A�֐z}�z�#l�_���	�C73�8�	��,:�A)R����6"��kA���LK��$
�3}L(�$i����E�Ȩ�%-en9L�C����>�1p񵇊�C��֥���S˱Y�{��o�mF1�R
N����D�Y�x�c ,D�wk�%H�����E��x�����<�:�v��e��q����G&��O���̿���C�~�~A����C��a�7n��,V�e#԰u:�1:R��wr|���y���J<v��;�<N�`���Rw��):B@?5&��2�ּ��*f�eN*q���ii%����/#�W�$B �P"9{�F��V�D��ؼx��·�e�:�G-��G|`���{!x�5�8OP��I�P��:9� 덎kƘ��1�ؔ���-LAn ��H6�~
[���%�(�7���y�����P��t�����,�|�2z�?������'�X�{D%NV�t�iUZ4�;�G@�|�f�m\҉=j(���Ө��C��^��	g�_� �!�u�.qa������}��al*�XTo#��S�9kՋ�+�?+p�>�{~	l�'0\N�ن8BJ��N�����;��.,e$)M+4��G��` �.�Z�4�r�!�a}�1�����+�Q*ag��`�U2��+k��d���
�����%Vi�Db�|i*7�@��"�nn'CႸ'#�o�jۂw�!�	;q`��GցKa�V��y�d`�΂�$*-q0�C���Gꈩd$]ɉ/J����J���q��[U>����������zIEz���i�F��l�rV�2=[na�rս+ىy!M��o��Ы9�q��n��� ��~����ح���fU�J��W��V���(�D�����Q��W�.ۻj%&N�޻�@����u�Q#�'1��e��?m��?~?��k7̈́Q(k: t:�q�:�
���J�^����e�����W�L����7L�`B�p��C�#�Ogo97{���%dv��8�^\NTm��q�Xלw�: ���KdP�S7�q/���ww�4?��'��{^f���*���y��*x��x��x��R�$A%�l,�6AJ�����/��s8w�ͯ�fۃ9m	v�(�B��q�q��rV����c�wiWÍ�"��13[�rj{���r(ol�5���Oc�V[,zT��Xd���"��R~]=���g��{%Zt]�a����K�s���<�~R��l-�xz
�7�\�+�:���zY>�pԙ�x�����`����������eF���x&LѢ�i�Q�l�fģF�y}"�7�9�e�짨(;�ǲ&��##I���^'y�T�"���)-�)����c�B�^5�1�;�,��l������x�v�%�!y�7\����8��ٹj	��y���1Ց�%#��z;�YU�@:���P���]��	�>A�����H���]#3G�N '� b�#��P�_,\����w��+M4΋�<�GZl�i����Y���d����ew#78�u>d3�(73X4�xU�:x?~I8�A)BڙQ6�%It,r�5�6�������N�z�Q%K���3��w�#t�B��5�߱Y���:�ܾ���\ç�l�E�"����;nAh��G�N�4��3hw��2#!6� �h��]����3�-^��|x^�3u�4ai��֒f�,f�^F��>��Ty�X
�P�;�=��W}Ѧ���D�яU�XT����=�a��X���a��ZYv�l5�.�Qo�S��^U�������D4>�Ѫ?=��������d�����>��R�3��72���&mUu22�kݯ��+*ffkZn_~��75�`ExkA�K�-�y��hB��'�0�[yVA�P�e��8lR�m ��Zڇ��4�K����?��ѱ��v���\,����c����Yw ��{����ep��������c7��))���ˡ�	�����9�g,��)P�Tgz���'��W%��d�A��dİϊ��k�ꓜ��1=�o_	|Yef���1=�`�y��3B���F~in����Ƥ>Z!{��'��R�ck��S �q"���8��s��#��l��&i1��~����Ƒ^^��O�'Vh �T@�� [M���f�mĢϙ(�>{]��Z�0��1�fn0a��\e��he�R7�z`ș�.���M��y���ڑzO]h[z����(ϑP�Q��D��֠��GO�{��2.��u/��!�L{>Ud�01U���n�ᏞٻyѬ֌�C�d�T'�h�vv�Rƃl���TS	a�!�9z'o��Ȩ���k���2͒���'��R6���m����X\3�>���X��-cl�����:�g�ԢoīϦ��:.�q��Fl���T8e�x��Z��Լ��C���Ĩ�i<�pL)�WM��Kհ��]'ݥ���m\�B1�x�a,���*�u�@��&�.(+�Un�HeFa��6V���v0�F:ltC ���9KYwJ��We��3��#R�$N5wa�gD�*f6+6%{E^B`�Z�C�'g�z/�wie��g5�A7zI���Њ�A)o.�K#;
ִ^��Ȃ�6d�޿�Ts�Sӊ�nT�I�R��D�e:�D�xO:��CA�`��}�3�2�bw���iJ�:K�O�mx%�ҩ(��X=�е�'=9`M�:�-\�f��n��q�w���s�(T�NQ�\rz@�,���#���KD���R؎J}q�y�0W/+Wѧ��P�^|���΁�����	3���۲���`s������/� M��Qx���ʇ�] (^��zk���	������9|O��)<XF��N��Q�	�6��0��tMI;XY����d+��q��d)+�Qq%�3��G�>��	����yx���8R��R��*^g�q	M�%tW ��qr��9C���Y3��������S�-�������@p�Sk�g�iC�Ma4�Z�xW�cS��4Jq�g�I��r�7�5'J��H%�$�3�o���&a�h#8����4:���rzq��:� :v��\O�ÔvR��E��A��h���#�`�,��2�"�F��������R�-c@p���ٚf|M�/�7K�@�yE��Y��lL�+���\��*��ٺ��3�A�N���d뭓U��̌���	��BD�)�0��p���\�tm.�:%Cd�~����e��ٚȊ�3>�_j��9?܊�?2��A$�:�����ۺE���菒�#w�|PoA��Ô��?Sȩ\�z��'I�*��7�џn��/�2��Ƥa�4�Ξ�W�i��o��n��ه�uM?��s��rָ
�9j��i���/���?MbA�aԤ֢��z�F�/_I��`_�If�-ͥ����@�����=�u{�ܾ9%���F���5o��Ywe9���gP���`�y�'�176�Krw��C��=ٵ���7�}���R�\=�;a�,&x/�q�A�]�W�Ja��C|}�/�A��R#6�{֥�A6m�߰0����M����9��dҰ�e?ϣ�����g?p��?�z'�S<k��q��eJ����#��x�E&�
JK����x��C�
��v9ĳz�d45��X	d{A�WÌF#��8D �����BU��r��z��"�Ք/&���\vrm��o����.#pG�c A���O7�y�f� /�G�����5M�N4�	f�����{1%WFx��t?�b�庩|�v�T��!��.g�NA���h���}�p�-�n�&��0��šX�E����Ǻ'a�.�^k�,�Y���ji�^f��U�[�t�����Z�#rg�9�7��g9�W��n�bG���D!��R॔B�����f�7��r���"wr��'�1�U�%�=���l/�f���E/1ɵ�|62��Y�ޡc�ֽ�\|��Ű��=�!�ֿ��Ƙ�9h5Ƽv�8:t���:0�]����k��R�d�������.���"�G��ΐ�zb���,�E�\��I�0��_r��=�S�� �� ����5�`�5W<��uj��cÞ�n�K�ڍu�?�W�$[�~��CӼ� a|=.d-/ofׄmL+�<'d ��M1�+u���vK>d��s�����KD�z��N�.�5;�3��8:��g��W�;���G���|�3�o"No-��Y�(O����{�#���E�&gʵs��ӕ�T�U>���*����"�E=Z0JƑ�;8�O|�w6�}�WN��(��[T�_�Q�pv��;��q���&~��i^v>�O54�2H�xݹ+�����F��}��$vj��qBL�jL,hl���J�l�w}ϰ�ղ*Dt_��]�Ƅ"�����]7�ߠ�`.����9lof+S8ٱ�y�M�Ս`��., jC�qE�	���/�6j�T��u��\�@����<o����UB޸$;z���3[@���a��;���Y�$`��$_�#�x�'�V�S=h�!�\��P�A�)��L��[ʿ�9d�.\��X����A}_�9��,";1 � ����d?�E�Em�͏G?�e�:k�j���2��M��K���d���d^6v�馎M
x$x�e���1�-�-����_�ڠer3�+��	v!��'-G�|��f�n��w<�B�c]����p�$��ߔ��0�Z�Ò_��n�d(� ��PzGK���B�r��!�"7`�QH��f!��0��s��^9	�����x�㓫V0{�ݜ�1Ĉ|f��YLÉ�P+��8�^B�n��3�P�����$�U�,3G�	I�m�O�ls7\0�H������(s�#�jlg�㣽��,��3�ˮ"�r$}�����GǪ����+�ݵ[���b��یCZ�����!BA�_��?.��T�&��I�2�d�'~"���F��B��ZRb�Q�2��ģ�T�oܶ�f��C�<jw�WZ��73�h�^2�a޲��g�A��������s~�F�lY�"�s��
����=����\����(���x�ʙ��'�\��z(	�n��2�Y�n	�c�^��8�43�p�p���	Q�J��Z��Sl�G�;�ؚ���E�T�T�b���ɜ�pi�L˲A�o���Ϻ?�(ˊ]�_-�,�S[�@~���A�z:�Q\�nk�;��!,�k��l�#�*����V����88z-�+y���M��A�6�
���X�`C@u�%*��B�¸��l�R��:}��ձe "���m�OU����5��Bjڏff�:N�D�'��X��xi
ޭ��M��q�}���_+O�����e֓�.�9���p��f��g��ୃ�:������'�{��m\�0�aYI8��z�#瞷�!�K���0��`N�GO���o�7Z��P��-a}�-p*J�颕�
�`�4��,	��
��k�-��@��ۍ�����M2M!�A����eb��KYt]��+��W���n�[��x**��$� ���WaQ�>]Χ�"�ש�+6�c���e��,�>�w�I�u�ݮ����#/�%g���*~��,g[�ȅ�aݵ+k����!t����e?\�#j�D�LJ�GK��2K9*��I�N��)��
%�S����2�طPM��+v����I�Շ�7��B��Z�o��<�2#Qjc�w�.��H���j2}_&��/�&��4��u_�h����N�����S;	<��۹M�E{�y}�6���[��ذo}E=W8��(�=Y6M�%z�mZn�����36�R�"2�H��MM5�w��t�C�^��/��ƹ;�pQ�x9�!Hb4����ʴGl$�ŒTߤ��0RE��H�\I�&7Y1��s��T')Z�Y���BD����>�B����7�o�9yj���e���-2��< �lOdwJf`H�˞�vu���.�n�_L$�J7:N�����|#�%���o7�ٕ�����M�%��!+����\EY�����IY��F�ݜJ�5�����gW�"?E��g�#�6���ݱS��$��'�y�$��7Ũ"�Xi���^��N�z�V6�������rE̫���Zr��'įQ���6>^4�� ��ajF��х-�qLӀe���I Rj="J��27�w�B�&l�L��w/@���M��.\4�����NSt!�b��玻�L��X�����5��D&��� ���X����l͹��͇�v�p�^ji��i����v5�.`��E᢭�x㩳����-3�5-�ǧ�r�� =�y��!���|)��T;��>�o[_vz�A�~�`�3_Skt����m�3g�s� �7��������7�"c;O�:���.p�V�,����ɶ�9&ch�����y�u�D3m%+jb���LD&Vrc�_RP�C."�
��&�X~��g'2_T�eL-~DY�֨*�9(�&@�zb�R���w�7C�wGj;qX�Y����Lg�xg���Y��X�6�+��N*���-4)Q
�ͻx�gY��Ґ��d_	�����٥��x�BceX�r$�3*�3+b�0���'jZa����fv,ek,ST���iX9!�Z1�����e*���f��w	�8�b|���^�2����\ܢ������7@�1ӣf��nb��'�Cd��g��,��*�r��L����K���kyR�^b+��V��k O�x�Dn-7` '�X�V��[9�>b���?�E�֩:ʁ?�dː�I�L��b{²��j]�9v�U8�R	+[U���3�Y�l��D�}���[���$�Ϊ�hWs����ԙ������A�� '�L����Ԍ'j��m=V�b��r {V˺�y��:΂���VAu�i}V`k{��!�c��_��I��m��V�`+XU���nb����wػ���	cL�ܪ��}19�`�V	��JXW�o�Y��Mg�Y�L���b�-��K�O�{	�p����pAۀF�,�#��D-�
�-OA����I�Ar����"lI��tz�:ޘM�	����8���	"1�;+	c�@����x��e+}<G�WX����܄SuD�h�Ӳ+V-�E/]�5^���p��3Z7��� ����R�G��}���m.�g��J��*�t��n�C�o@CP͆�� �Y�G>�ŏ���x�a=�x:͡<b�=��I�a-�i���Y���>s��!�BU匁f��7)榗@�NA�03��֌v���"5�w?@�ªՅd���R���5�f��5z6�g�+���|���{���>�B^,�ܽp����&"Q1�|b�]d�t�6U�y�v	rm�b��̎�[;ew9̨��U���OQL���� �#<��w�����[�������Z'=�z�i@�˃�	hs�D.h�~��OU�ߟ�������s�B���O%�8�pNB��Ʈ�]��~�i����C7�9��&5�;D��;�E����� ;�7�=W>��Vz�Zx�  ǅ�z��Tޟ*~[�U�m�w*��B���g[9h|zqD��T�'��Ӫu��|47~ÃPM��z��o�>��^�U4�C?t���h�E�R��
s�ՕO���"�d�'~C��d}k���l@�������������T6����c��9؇���Q�)g�;�Ek\�#�3^H�
�Pd�� ������X����9��k%�{u�E�y����$�elw��Ǳ�	a�c�[ą��'3���7����G�T�[��I� �-X�&�AU F��O���4WY�l$. �]��0	�ľ��c�'8���
�����~�=YI&J�#1m2��}&d��}�۱@�ߘ�.M�IQ�V�٣����tjj3^�ט(���t��DX��J��|�6�M��'��)!�o���ݑ �������
�n�U%��;��,3� ��=�E���tZ,��)/�/E��R*���:�΁�������>b�nǖ�Y��*^zb<EX���Lj-Q_�Pm��4o5�%m��g`�|=j�{���~�3��sh� X�*�׺�'{�s%�^G/�Kd�p�;bh�N�6�����,�9��Rc���B��K��`�F- ���%J���+YO�;_ԪG�0�^���M�=}AT���q	�Lԧ^o��+�Vg�d�Wv��9;3<�O(�f_�h4R٥�$MI�f���:	
�pKL�V�:�#��"v����iO�A�lxjd�t��IA}3Af<:|g����VR9(C�������Z���,Ŷt�>��~+s1�I�O��G-CX�"ۘv�����C�)��MUDG��ѩ�Ϡ)TE�ݖ\%dw̑����Nܲ��0ze�SX�Z�O~L/�Ϲ�8���j�_/���nF�h�YNY��QT$�1c� 꺶��g�פ��=7~�0C�D�w�b�?���껇y�����y����+qn[��9�?�"�>���OɄO�O�n*�f�YP�C��?Zv�>{\�e��r�� �X�$�nl_ğ����g[b��L?e_��ҩ�D�ܸ��L�=�V�T��k
�/<���so��Nw�p���굑��A0�>"4� ��T�<��G㱅"Ny��ʟ*v:+���0���L����<^3���"y,N�.Iu����x��r���8S~Q�����y��˙?	(��ېk,�8jՁ^@��j�&���(��x���'Y�	P9D58]fL�20���B�0���Z/Hl*F�)a|<��L�.,��ǳk)4Se\*q�X5飄ˌ�&���)��w�v��ܟ3θWŭ���|�:���qF�,�t��;B�R0�i~��sH��]"B�\���@Íf3rO	�����1�/���OW����>BX4V.�����z[J�t5��;t���`6,�G�w☙#�NRǋ���c��l�s��hο�lLkK \��&-���͠u?|�pC-���i�9T���;��ҫ{gO5	����`���Ȭns�Gш��6zm`Z&�!2�g��i�q`\z��&�kZQc^�#�f�{����
Ek�DO��i>@aq����1�6�&��Ť�d�"`�G��#L�k�޺�SeC�x7:� h�$�3��Ol�`b?�$y؅���YB�#<�e_`Ϻ�x4��u��*�����]�[�F�&Y��l"R����t��E�����Zƀ�s��H^��H29p��Ł�E#1��)s��t�ե����W�SV�/v�$2t"�L@Þ�A/�U�y	�v7%n�@
N�fz�KU�Pg�_3O�^Я�΋��B�m#�E�n��������%X���d����!3���أ�ᛤc��0���C�,��`%���g��A����2�(&�󷖿�gIW���C��x8��ea���K_E&O�í5��;�p�����X�U��`_#�I)��?���r���GM�B�K�A��L+i�̏)��c��\[�(h�<���"j�s�5~LUB��Т�c��P��i�����J���:���$K+��S�>�#�K��>�?G+m��s�Z;�V�N��wl��xMT{���.n<�'��`#�j��P[���~D���ó������h�k1�<�*l���:�j��K�/a ߔ�z_���G��-
��*kg�q�z?Ϛ^ARQ?�%�ݙ|	�z(����%a��_�ed��z	/�쐆�)'o:h�u!W���ж�0�Kp�zkE��|A����q��>���~=Υ5�uR4�Q��b���K+�.9S��nGn~�؂��S��"�j3yr��p�l�&�>�=a_��S��^>���#�Ǉi��d��;L��]��,���;_�*Y��-�V%���:�o"��U����*��-�X!�����%���~�}�eθ=�f��ƫ!�o��R�>�
�g��ܨIO �҆�/��W_Sm��]��8�\������(�@|{�L���hq��P��{cR`f\c�9	�k\70yI+m�lA�/�Y���`��_��uEt����M����/�O���$=��{�jw]�74ou��h��ښ|��IY'|+�#�~�n&ݷZ�:=6����lcg{���3f�5�O�ざ$��Q!�4{S��ڥ��e[��	N�Ou������q/�dnLi� ��+�8ת��L=����>�N��ze5�[pѤ�g�+���]-a0�ɖܱ���AO+JS���xS����C��_��נ�5���N[���W�����������Kw��<艩��X�8�
9��hxs�����̏��������W&*�c��CU#-��6��1��e���Ck�_�jb���7 ?s��%�b�A?�0�?2��
S��+��VA�ȼ���kw��	 �'��k!o�k)�,���@�7��<k��O����4/#����`�Pg��|�Ή����f��d>�U�~� er�e1�yN1�t�w0���b>����;�,�c��I�ڭ��]��dhC�1h�7��T�LO��&Y��;������� �D��3�A]���8U;��8̲ ��x�!�*kw�oxr+�l��u�����'GOW�����0����Z��9�����T�w�	�l��Rc#�g��hG�9�Z�#�:oN��Us�}�:��D8@�j.�����;���_�H3�;�����uA�
-˵��3tai0����xM&�S�P���_Q�����Fj��p�4sSO�IX���Ad�,K�������2�sI���/� �c�v�����R��<��	��g[��Xj������K���MRP)C �x��[��O�F��� r�	���4,!�/A��C0��w�	�^qpTT���h{6��RJ^	�,����Ѳ��&���a�UB�y%��ѫ;�wUݺ�Ʃ��le� ⪝H�K3Fį:^�v�\4M�3>�s�Q��%uбU�r@\��K��aE�vץ�T�.B��4�����ߴ�]��r��Rd�%
��N8 �qX�1y{���^��n9z"-�3*�qڸ,�y�����pѕ���*Z��81��e�*N�=�M�[���׌
��-�d���3[�n�;Z��m�kKG�H0E뉾T�7ũ�v�����\k�Lt�5��D;��f�
6ۏ�+�58#:���r*��+X�4�A����L	��M��2��6�,�aL����6zˋ�0O���v��.f�L�K����a���/�(���8PH��%����o� O�т]��צ�1R%��)�3{�p�J���+w�����!ʱZsJKz��V%ES�pM�I��r�=Fj�b��ߥ)4����*I͎��o_8@i�{��׸�{A�:�csx���;3$����)8Q:��R��	��C1��~rډw����;�iB��^� ������7�v���Tw+5r���P�h/:��\CS<sr��i��e-˵�v�¤�ƫ"aR��$�[߷_Y�Y����HW�~d�Z��d�U��tF>4l���^�ʨy,Ԍ�g,$	穱�QK��*]���-�!��y�/R����	�\P�5���zs�]�aH{�O�&��y-�!*��T`�^��8~y�Q.u߉ȯv�*��6�鄋4�䚶
)�{��Z3j�:���gb)��-�)��|��M���U��qXJ���,�ŧ��,�0�u����kP������V���e�Q$���ɖ:�|�ǚW����Γ��I���sb��r`��sy{��K�; LRF6����`ye���˥�YW�3�ϵX|��-څ͠R��х��׍�����R�h�hu�7��I7�֛`S3�u�3�$�0c���s��|���Mx��}�	n�m �>���Y��1*����	'}<�P
�צ.}=Y����+ c w}C�H�O|q��"�wr!�F�RE�$�E�D��ρ�^U|tG�p�����%h��
K�h|֊�M!�w�n������X�JB+���*��I���!�y�/?��'n�).�(p��z�Ӄ�︨|��3e�f�������t���Y��C[8�9��T��&�=�ǧ]��EA���Փ5�����:Q��<)�t�̪3M�u���nr<茍d��i9K�ٻn�G�vn��LD̓�S�TM8� 7�D_g;k����m��gྰ�8���;�[9�{F����;l7]�����i��vf�x�h������J�"o��!�&���,���"}�T���H1<����lV��(S��@*�֦�dE�����b�m�\;Y.Ha���$j2����z��a�a�'�����˖�\����a�wn����ͽ����"��
�D��ibOX{Z�P�����5m��Bo����p`�iV[�)m�y'��Ȉ��@�}D:ys�#�g��ռl�A1r�a%Q�d���G�����>�υ40���2�ϳ�}���&�����P?���b r94Y;�zy��	~�$��Zk�|���(Z��sR�9���D~��p���4s4�0�qJy�Cgjd�1�C-3: �~���KC�hHB
,c]p�%�3H^��ƐT�=w�/A��?��rL��$�)�d��"!t���i5Oҝp.:�JY��Pc�Y���RI#�J^�x��'�X��A�I�Z@��M�g���W�U����*��/=`��Ժ �K�i�Q�����.�( ��n=s�,�u�C�f�t�
�W#@����(�3��el,�.�D��!![���n�~��QW{�;涟�� }���$˲F��Ks
��o	��(I7&	�I���|[4��a�~�>V���)u�:�H�傍���5�@�#hU����j-��Kx�Ʈ:Ѥ����mR]������|��.�I*�A����(� �6��D��.o���+rKr���MaX�ssM|��;H�1��h���N3;�����}�7�->~�?�Dң3�-xt5�"�К�����<c9!��L�Q�KN<}-/�<=�҈R@�t������X	+I
*�Gv	��W1�lp8�oK�KK��7���WF؀�躎!���d9���"��x}�־��^j�MF ��-^�}����G�>�l���B���ӯU��*<����GT8<�o����.���|%�xl� �:��n�xA�/�{��/$�L�����w�2G��*��f��qJ�6�d�
���Z=R:�Ҥl�P@Cʗ�48�2�0CiJ��#&�<�vm`l���8��E�~a9�q�[ �҅�r16ED��B��c�Eݽ�
�"J���0���K�4���ұ#y*Ђ��Hq����[i	��L�q�:��
���_�Z &�1�Iȑ�T�ŒF����%%�^�4�p4�^��~���� h���j_h뉸��U����7�؁/tJXy���j�z��U�WC<,�N!QJ��`+XP߷8ocM���9��w���QV��*r(��f�}6�HL���I~���a-|�F+O@�'؛�\���j+������:e/O�k��S��
�������:����ܣ/ҘZe��,�����%,��/*�o�+	%��A�ߤ1b�5E��%OH�Pr|M1N��J������D+�\%���h�ߒy�7�g͍���<��&OU>?X��o'����WSa#�ɛ]�����Qز���b�P� � M�i�-�H�+0�ِ��{�Q�3��^�\��}�F�f�[�0V��/�"�V>7���zqt�|��\�`a_������M�j\]����J�r[*[���E'^"v�����47m{G�۹JO���y����w��hp�:S傦�{Q�k�y837�AEK�3yƆ�%Zw��i}�%��At��<�_J5��g�M�^�X���\m?�1���?`�� ���n|����&��\{K���'����-�l v�i��c�ܠcA����f;U�D@F+��㏁f�n	��Շ�w��YXO^��`��o��bB������亱4��1��L#T�Q��|���t����z�ޠxi�q��@8��?a�S$uxQ�V�������|�6M>�٘85a�3��:ף�>�>Xb(#�Ȗ����9:)N����	����9j�Ѷ�|�,�"��A�,��H���ڊ����w���eL#m��Fn�ҵ��O�[r�j� �j����q��c�<a�Y��0Y��
�w��fT��iL��i�h�ې[�\�����ek���.�����]2�*���X���H��ύs�I��R� P��zW�kz�Kac' ��|oX\������a	2�Y�o�^��1���S}5]b�m��s���F�?��[Z�)Z�_�>�h�=�35�]D���6�Չ�ɠ����L�a���c��B�Yx����3Z�����8vr��c������[�܆KNƺڶ�W�^�&����P�[u���I�K�(�p���W��9ޣ�������e��{�kW�R�Ao+r5}���W���R��,����[#'	�}�,܄��� ���u�eJ��&Á��?��A��Wr�:�e%�2#]����k����ͪ�ȡ��;p_~V}/�����w�t�	+=3�%`<7Q�G�!�s��_|q�+ѱ��V������f��/�=ګG�=���x�2½xm��S{��'8Pi3o20��	�������R�/�1��0���d¯��w~���62N��d~\��HMH��,?���6(<R�����(���p��l/sh��|��ɓϽ����#.��ʻ�X���}���I�YʖĄ��ҝ���� Y*��%n���#z01�9�N.�C�L�NE`��E�p�9�P!����F�d� �L�Z�8�S|�v 1�����lƤ#��z�N+*��#���P�$���S��Bt��e��)��-�s��w�tH�)�L+��nug�}����a����X�Ϣ�!�rf���9K�V�wj8��Y$��9_� �1����a/��x��ts@�K�AyO�k%�6���C���@�=�̖KM�^?�W���Hȱ���Ռ�.�.���i�,�/=ɅnW?y�$ۓ��_@�:Ե���J#]�|��I�T�@��w,Mb�O��b��c�{Li������
�	�b�MH"y���gǳ!�����F����-*�[�Q�����=� �}��~����a�oJKQ�b��.Z�{���&�v��5Uܱ���s��LL���8Į�s|P��"�듬X@]�""3x3��s�k;A뀋�Ҋ�)?! ����2eMu{c���eY���J�h�nK�6�Nl�Zp��!Vh�Z�|#����l+����|�0�
b�s����*��$�o�� ��ڒ��5���)'Ұ<�_�L{�,���M	
�/RrN|�n��Rc��fIVa�K�/F���:C�KD4\�=/SB�zm��3�L�Z����s�ɨE*[{��FxgG&�0�mO3~��>����,�tc3w|�Y��or���DHO��x���}*8"�$�3i!8 ���L��6c[��,L���~�G��~	�HL�:��!� F���mi��~�Y{�T�ͱ�R&s>�؜�D�s��(g����ԉy�5Xl�s�����y�!yk/�ƐPk&'0w���b�ۡ��O�}|�se~.	%����]踘�5=z-i.� �.����)a
9�\jL�G=Hu���n�Wd�Q��ڪ=f�mź�����j1B-vƌ[���bX�Q�N�g�*A�o5gs����`��Nl�����6(ɨ��@H��y} ���V�k�if��n�!��(��v��S�Sd!�Y�#ɻ��.�C��0���Ը��#[�X$vw�W��toG ��Ik��:Q|yWL�ʱ}�F�MH�v�[RZ�>4�W��a�~"�}��U`p��&�G��׷�[��f�&)2̋�xM]fD7�� �S�&,�l���gR'*h;�:W�MA����D=(.$�-+�p�~���x�y	�5���~��[хW�� I��tW_�u���. ?����*�۬ D�Q`������P���W�<���"9w�t�� ��� ��s������gW Xy0��'�Fxk4�������FnI���m؟f�[/��"^#b,N�Е�f��t�A�O�s�M�0�<?NJ�x�N;P�n`N$�ڦ�@}#�a��Li_�O��e��L�j�s�]o�c��u��P=y"��)��JZ����j��2(��$�c;�����8�"�u��q��� @T:u}&Q���}��5U�%[� �O�!5�����+���k���T�K���1�w�OGJ�X=(RB��6��e�����"���^2բy�@��[�f�:d��-r�jiWV�c-9qn�hg RU�n�Trk��Oj�%N��Y�i_4ͤl	�3�C-�Ʈ1�$��_sW�V��m�[<<T�ր]��A�1 ��&���JX�;0��œ�;������~j�G�m�(X{sɚ��u��g�F�h	�t��-ݑA�R�d|�a��T��Uj�"�b��ȃ���B��"�.��PL�P������?߬�����ȞM���j��/ͷ�J�]œ�!�E��Yh`m7���f���_'Q=����� 1���}�&Ȁ�%ݼ�N��e�<���� ��dE�MY������%�I� )!�Y���=�3^:�{^E]g��NưK�(������zJ��.�������iZ���-��HZf��G � ���d�~�ln"e�����y4oe���6�t[Y����������z�'�@�?�|�Z����Ԥ<㳓��s_g�����'숷�_�6�P5�\]g�D���u@n/"$%����`�i����@��B����T��0��M*�.>f=���~����KA��6x���M��c�=/��c�ϭz�	O>��m@i�M�e8.����NӠ撐:��V������>�~x3r�mS|+��ޙ=%�٫�?���3�@V��i���z:>�]H�V���\��>T,j?{G�I,�_oa�����cp"��^O Zw��:�<��;۠�ٍ���r�~�����8D��&��>�֋��>�@�JV�ф �r��֧�b�4��!���/ �n�ϳ�{2������5B�����b��5	{{��+ū�kyI���'_�g8?�U�ʗ>�5#-/��|#��i�I�a��c�
�Þ3
;��5��毖=����n�� ���@�%�RZm�۬V�G"�fD�Ez���jnK��Hd�;�/����m�|�<��<	��|VL/�`�q�Ԡ!쓹�1vi�&Zs-pɸ��CoQ�n���=�[kF���hz]�����;�i�)�F��
�#�i����?�YG�0)!������m <�|��\sJ�FYXs�Z�yz����P%�� v�m�+�D_Ƽ@�ˤJ��Uf�A��9���;��z����l�ª����\����;�@�FJ=�/�����ʏ��Z�YS�/�&���ʮ�	-A}������7���	Z� -Hɦ���)Pn�IQ�t#h�V�tM��#,=�q���cT(���k|�!{E7����E��ufI��<FԦ�#}"q,mڅ���n�o��5YD^��� �g9�b/�)����B���j�_��,�k��$x*��,�:oQ��;Mǚ�󍩦����ڵn2J��M���7��YkI"�ߌ������^���_&'��4�^�S�خ��-��߮�6竑��.;qL=�י���f�X�;�>@7��e\� o�|����V���#��&j��.?��aW��y>�00�ǻȏb�Ol�j�3ȳP� P0��	�a	PB�
d'����b���$����(�g���Yr����S�`�n�������?�؝�WP����'�w �2.�Zxr>�+ۙ���V\���}�Pql�F�ڼ�f����F[�ƅ�|JP�y�KA0�lE�hJE{�AP�2
>��� �+�9^��=��$����*���!)|��)���(i;~�����ϭ&���o�e�Q�b�]����e�\w� P�ꤺ�u��y����}$��(Op�):4���+��p<*��E�F�� �!)�cغv��b�w��Z��R�>��`��w2b&UBw^�}�ZV��^T*Dfֳ���+m��~��2��%G�#O�-��]GLA<y�e�V��V�S�{H�ZD��^�<�`�<ƌ�=l����ݫٱ�5���Zd���Dwq�Q	_f ���8�Ⰾ*,�*`[�u�C��ߏ>���W��_��pI��x����*~pʯ'��xR�Xh�����iË����$-�2�R9���P΄(�J�b�u�LD[J����ȑ	�+�(8T�r�8���(Ae���&��� zC�e10�Q�3���І�N��wq1���@[��>N�0
�$������T�����`=�r����\~�{���`��%�������.#nyt4Xx0��!��6�獹T }v�������m��"�����fe�%}�����9�jm��$8m�l��Bd�ibh� 8��x�[Ϳ�ՁWv3#f��4�>?Xw�`��a�vR�o���SP
�����%Z�x�^�
��^h7C�hk�˴�ɋ��D�E��"�H�I"0��U� r//%@{�J��� �ߑm���ڤ���-Ȯ��D?��T���,��{I���v�쥹�HP���h�vJ�����>�L�q��$���؇�75g�>�V�D-�vIi켄��d�$�Z9
�'�Q7��Nk-5�a�`�%�:��!�jʰ���-1���
��Ԯ�r�NM�M�gk��~���Pz*J�b�5��"_���5Lp'x��+�G��O�Z�b�Z��PX��l%t+H��`\1�"Ur,U�f��2U��,ȍVx�	�%�N�
�r/����}E�'�*�i�ޖ�,$A[$h4�1�s\:�����F)�U�ߡ�ڕǉ5W����ā2��@x�:��JV���@Ӂ��|=~����%�:s�m��]X�*)&�`��5f|��jg}�]�dr�����-Q��h���s�Ϭ۽����	LLx%h]Ђ�x�l~�畊A矼��V�H��%0��/�AOji��?�p�y�;�D��s6UO@,�B[x0q�O�s
�{�8���b>_hQh�����|3�]���ץ�Q�Y����If%�#�j���y�r�9����(7%c�)��ӆpB6S7�[�憴$�	�����ϒߡo½�X�*~\7���?^{krMC�BYzq;���'�����&������G0�-){:p�*���]&���S,iJ��J>p�q.���@�Y�}���-���Z��p��������o7`(��1�p�^�owr�$�4K��E�����\1�t.�z���C��"&&;�h�3k��@֟�P�:����wV��v�"��ux�n]���s]!+��:���S"���V΃jI���;C�F�Vuz��G7c��k�a��� 7捸}(|�|'PN˷7��C������um �R��F[�;�BYp������s��l�YJ��e�w�ݧB`�L��#̽�^�ݝj�M����`��Í'���iUA����5-�T³�oo{�Ł��%���������6C"�1}M���4��Jۚ�+r�p7�
4��b�\G`�j��n�����x��7�5@���SA�Tkj"��[�2�~��f��dh/r������|n����w���Sa��Os3���̞~Ջ������ۼIjo.�CA����� �ј^�)��q��ǿ��r����j��9� |�@��;ź�M�T	ë�
Z;�nJY��V��L2�n���v� K��:̲+����fj����mU�M��������fZ�4��XS���԰���:~�x67	_�(jpHf<{�!��S�QC�_]޸��Z�N6�
�B{�������<����@��vwD��6���/���2��j�e���������!�\�L�a�����k~M4�g��\���t��T[n[�6�q�!ǝ��h�!�q�C�q� -�e)��AQ�� Ƭ-c����	�$�gh���\,����p9Wi������vP���'�����	�L���n2H�7��9�V���&���K�!h[��zƭ��-^����4ҳ/K�Ƀ&�"��lH�G|*������{eЙ���
$=�>7g����S��u��ӑ��
��1Q�*Vp�t8Wɗ��U��IZ��`�/ن:n�{��T�r��3�mO;���4�y�8땽��c�x��B�0s��W�>y������I��f��F����b���Qb+�(��"
'kM��JF6z@��-��Q����Պ�
&���\&��}�
.\"KvaT�gRS4�&N�pX�.���ܶ�>Z@��,%g��r,�4amEQ�!� V��_&����g���P��U�W�c!�_D����)d]��KHQ^}Ãz�u�K�����\C�	��������w*b|YǄ �.��ĭ��.]�7�
S�{���u���/�e�.R�-���}�������T�3rɬ��=�,��
�Xh����j0�]3�r�񵝽A�'v�>[!˱j֭.th��'�����1�/�z�>���,5)O�w�9����.ժ�V;0�m9���n�M��&���x������ʸFm�W��*(XS�_�������u1�OU�pd���^"�Q/-��^N�#�¿6���z�m�ԍd!~���z'��$��E;��3�@�.���p���(|�%�,T��n���)����Z��L:J���')����s�>M]���>�i<�7�(lPU����fKc�V��-M�X]�Ix* ��U��aor:]Ӭ���Ru�C���c7��M��L�Z*��_\��.����zwVD̦d��D�q��:��+�Qr��k�:���~g���o�H����w�R6=GΞtE^��G���̙|��<�k��$��ti/����dԅ�a��O���JF}��S���ϛ�3���l�0��Ǉ��k|AB� +x�=!y�v,��+)lQO(��h/XKHB��Ee�[dc���	5�"����Ǔ0FN"�ޗ�N.L�G�틔��V^�5 ��1��d72m�uBfv���r�f[{AY�gi/���0��g5�{vUt����X���(��Pjȕ����Q�[����Z�w��c�)h�'�1�	��.g���~=
���iY8��]S�R��C.4��w��
����ۅ�kN~J����e��������w�Au��G
13"�)\ҫ�6f��ҿ[1	ħ+�P��/9!�Y��S�Ǯd�}�b��|���샿�C[��*���lٛ.\BO#n���ar�|���t	�T��a���e�F��4$f���+�@��� ���NJ�:���/�U����8�{�?2�z0�R�K�3G��CR����JDiD50�*��Q����w5 �R�F�����&̍�V*�^O�����(]|]R�;�P��^��yx�ݏ��\�^���!,䪋<�l M�,L��.�R���m�V�S��L���&%xY:��;i@���O��G@�4�����9���ս�C��
J���\��6� �E�G����V.��`���=���X��<�t�~#���-�z�NjO�!���6�B�6��߳��������|9���� =+ge�����O���d[�C%M#Ì�V.gp��V�yIv�2�i��Uk&�;kWx�uF��n�J}fG��:�ռ*��O����H��@� ��v&|�ɷ����W%�"E��*T�D�sGi.{'r�S�bq��ͼ��aX��c�E]��w�T��5\���m���0�e0#�:Y�^�ٞ;C�f��pS ���f��c]��9�<�	���/��-�d�!������~�-�.�;��M��]N����)�c�Y�з�V44-4=�)�;�"e��j���Rw}&.����j=�l��)��M���*��:���HsyY�H�yu�ͷu��j���P
=s�aD���w�9e����G������S�+>2'�3�H��E����.���q2�2pɄDQG�R-쐬�0���2(�����OR��V�˂�[	^L6����^��̅��p��u�)m١��v�����C���;%��ؗ��]����/��}�Nn���o�YtZ*S�x۹�8[����n9���raV:f�Q��p^G6}��NX��KB��-��d���:�Gf2M<��Ss�^�;�f�!]5&��!e_9�l|�g�����<�qy�/��zm�c��	��6��BB�hv�!|Q1#�=�(��2�L��zx��£ɾh��n��o)Q���{��3G�.z����%;�J�[w�ӻ�^p��<XS��EtCWuF��~�Q�b&�
jY�PUJIT��T�s�YϦBt��S��3,АB�?� �H���7��- �M�������<E� ;�DoQg��6����uJjJ���<o��;��6��2֯~���;ZX
��@�x8��V��j:�w�����㷎�H8�W��C�A��
H�n25�9UӬ���Pn�";��H2Nצ�˫%��wQ"�J��MXˁ�SK��*�9d��qB���k���/�t(kA৺}�-c��*�<�q�s�H��	��:#���6fښ�O�xv�W���q�D(��7
R� HdO3�$txߠ9 P5`����L(�2� '�����d��S�=���L<����7)4.	ۤt��:a��_�Ȏ��T
�Zj{M}<�}�������n�Qק�Υ(3=a�+Y��{�J��qgl�hF��#	>�~�N�>#�e!O>#,���_ ����2'{����|�;��`�>�,��0��3�R3��;�E�&b|]����<�~��ht���瀇�ws0q��o �N2��t��F��*V����ZM���f�B[�*)
͋&}�@�-��Hf꼵�a�G(-��J
�*�P�uG�q�C�z|�F<y�i\��(�D��d%C�KB��U�j���~�p����a���Z������e��aż�ܦ0��)lc��a%Ƈ�V�k�韕2e�l"
��A�����_�}�r���@zu�Q�]l��ݑ��=����2{xE�_����� ��(��Ln&�H#��F>��C�𧃬Ix �Q�a7�a�V"��7Ġ���mFy�_P���{�ZfJR�_T��a�pgUY˄���
w�޳B�������vw3�m���lov�� c��"��?���`B���X,3��}�i�F�8���M!Z#�f�2e��,k~X��kG�q�Ǭ���l�z��;�Zmu.���k�_�����`sS>�ŭw|���?yF�zd����S2�\i��d�87�c{�oj%f��$�L�l��[�R�̛��y�4R�-p8����ri�<�qP�F f?����Ǔ��k�@ǎld�w�\�w-WA>;����f��}![��{_��Vw��Êz����E���<`d�S�@�2��3@J�KH�ޒbW�L���~��;��7C&z�Y��Qfk�l��d�ޛ�ܠۼ�r��/��_\.օ�S�vn�i��֞�Bܘb�P 6X�a��i�c�mI�~㡘N�N���U\	
��ur��)�/�_��ή���V�P&QV1x��.4�"�i�1��%.1WA$��CQ�HU����:�ZH���*�@���;�+#��>v���$�w�o� �Ǩ$�j\O����w�
��h��W��F�T3�c�~w�w�����>
��Tn
��od�v�k,�=���l�y��7��|W�DT�+(�&/�G�KV�-�v^��,:��}�d�a�tY�Qa�	N�_�g ���HP!� @).5�Xwr��*K�5������.�73���C�J�T�ga�߿���n��Okc9��9��})�����~R�U�Y쉐ա�ί����X�@�J���ɫ��׎�*�<��'�����oǌ,lu��u�}mc/9�?�g����뇇�g�sj����pggV��hn��$_�)�����oS��\F1R��Ɍ�0�J�wFAt�.�P��%�J�;Am�=�M�,�7K�]">��w�Ɣ'���ඕO��P�x�db�m���FO�	LFP0��M�E��8��IF�O��6��R��NH���1�x�{����E��$�����s�����K�j��#p��鉈�V�7���E|lR�w�vo�����Y�h�6o0����6�dy��o�vGf�lu8��濕�Y�G\@�t��*a0L�=�k�V9��v&�"Kv��>���)�˫�[9���ck��ܦǪKe�x�@��I��2�������|E4��R���ﵲW�Zۤ���O1+�7��"o��u����k���l4uX�~Ǟ��З��V������]KkL2״�=��X#a��������gJնp��l �=_��,"f�f.RJr�A��#&܎����:QGnz�����\�ʅ����%%��D��M�U��+E$#2�8�3�Y*�sX���jr�	��me�Rȥ�W�V��H��{�"/�z��MVV��&��M?�T�-���'t<��V	�uN��^���Z��=�+յ2p�N!Ps�,o�/�̴���hE��Fk�a7�!�F���W�=c�y�1��}���i��Q�T�xǡ���
of�pe1����UԌ`��?+3`�̰�9u�%6�'<�m/Ǌ`[����9
����9E�j��zQ:'ͱj���X�A� �J����D&���s���8�aj��*6�y����b�8�Oŷh5<}i�3��]j��;���l�C��'�����L�HΫ��ٔ��}�}�i�u�w�Ǔ��j5*f��ζ�-uA�^�g��hroJ ��0�:�#4n�����'Hn�v�`���i�&i�EC�o��Ic5vE����7&�q�dB	7���6� ��P%�]��$>C��eNWHR�B�fJKpF���
N���42��5n���g��W�N!���N�)GI�����t���������|�C�;�!9"�Ħ_lDl\�d|i�[�h�#P_�������:�t[�ѿ���B�&j��YJ�(��i�F���[���R�R��Eb��˓��v&=:�� �adw�;���H�Vu���3.�o�P��ҧ�������RYR��aI;&g�%�r�� )Ȳ�{D��Ki��* Z>��5._�F>?�ٱ���
����Z8��^[���Ã�6ѼEYi�#=
%��;�WH
F�#V��c�Yw��uՄ|�a�H_� D�車�����c�\��"�_�=��p�*��Y��H���j��G|�o=[�w���u&��h�dL���<�n4}k!JϺ潺�!Y�yY�*�
ЀHUY�Y�0�r^�z�Z��ZΌ�	L[����DL<����q����dt@RT��@��N�����Φ.��T��͙����m���,;�+	��0i[ݭ��<*�^9�s�_��N.$Qvj+��G�<bR�G�$�����-�v��}�l�${�ʓS� �ٲ�Q��i��H�u7�3ɽ��)�n��D���W	y`�"�3��+�����'�1����{��tK��Լꃕd���^��jXRf�������cyW�B�ǰ�ҁ�T���f�֔�I]�����	���l�p��!+׹�&�m����ΈV�Lu��� ���br��\0`�
����ߟ[�#_8���lh�Ľ/C8�)������&ɶ�Z2��/���7I�]F���typˑV�v����@���1��^5��G�C}4u�qk�w��"��X�Y>D�S��wJ"<rx��!�X�T����L�3������j--��O���/)ff#�b�A�'�ƒ�ڹ�MEV3�i���I�3
G,��M3p�HY�mqJj�`�%�~m��k�
Č�������p�ت�) �T�T(Ԯ����4�ۂ��Lc��E� ���b/9��Eʵ��LH�a���Bz5P0��x��çQI�o�,���K�4�����G0/d���H�r�Y��*��"C̼"�����1�'�1_=��0�f�)������q���T���H�dˑ��d�s	lםq7 5&G[�^����㻷��@/nN���y�>]7��ɟ|[��9di�l0%�,���K�������V9*�v꼌3꥞�G(�$P����Z�z|-5fN��|(���Am&Mqi޴߉�EVtN
�@�~=��^��9�3�4��>w��Q�B�����`W11�:���_��K�s�O��j���o�Zȅ\�D�uL����)� >�	��|.M��Q� �7֧���l菺1	>���8�VW&>g��i��Ј����8���lk{�n�"%%$&��yG��c����
�ب��L,�)s�Z �?컣����r��e�Vis:R�4������g(p6)��s_�]�j��'�_��#	��Fm&�r��i����L&cC�@Is�O��)��,@����ǄJpe�03��?�G�,�h� �L!_FfRW�F���0��yM��0Ptx�&_ BO@Ë�W�f���1%8u%C)������)5O�n#\y��M�hN���b�8��*������9z2���Φ��F�t�,��ܺ},�8�
aM05�EԺ�O�����.�M�J@_�}\,��5j�&���c-�em (�<[��!ޏ�܃�>�a��]V�LM��`���0n�����sG+�L�?�KO��Qצ� ����0n]L1�!�#���B("�� ��a�`d�(m$
8����)�0J��H���?3R�7_����R��R����,6�:�2�� eb��?��gW�������1����	���� a3�@�%�@��w��Z	IEU�l�Q���*�V�2�����N_��Ac��h
��p�O���*i���6�N�:��`���Tx��9N��w�6�*�)�&�}e��J�J��9��	T�*I�2�e5�.@6�"e�@FT������[B����	��fa�d���&>����'�~8�>k��T+�"~�;���� ��%!isFV�|�P����RT���zg��V��$^Z�N�,���w�a��,4s���2�1[2�e����3��3�J��N�Gع�,a���mA�2�7׀�ھ*a���y'�=h��=��D�Q��q���n�ɏ%2���l�"�������%b{b�g���Z��g�����O��YC���;�Ț;*,c�3�q�O�������`��Wכ��$Ƅ�>tcX�	>��EX� ��ٌM��ޅ��ܼ�{�9��t�kr�ǧ�|��STT��� Y
���(�7Q~�]�c#,d�Rӎ�I~����z�9F����q#D#6{�c@[���;�A�u��žr��&�L������*ti�B�ڃPE���'�,��o�Ԍ�����ȣ�T4�o}�"�O�t��1�W���Hwy���v`ɺ$j�⪘zb8?���u��T���Z#}H]��MMx�g�,ݪ�uV��<ز{"E[��z���
]�2}��V,�ba9�g�I����1��#��aĭW�%�R��fvq<�àv���R����R�+���.�}�7K�T0�2��Ke�L���G	Do_�d�Ǩ`�7O��	&,��A��q�&�;�fF�]����������k�4tꥍӰ/�U���Z;	/QLq��eC�\�>y�-�q�ޭqQ��No���f�<�����O@3~��"Le�
/��-��2kU��%߯���In����>0Ց��/��xD- L3k6����*��$�6(�՟���aC�&B��'�Ė���+���'3�-�wPà�3�a~���}��["�#<>$?��PA�+�Y<!�-�w@�����!}[�ԀcI�l ��T���W��W��������n���2|p�[{��rK��s��D2�ǡ$�.z��W�k�^��qA��<���0B�K���!䓵E��G�ׯ��������A�1���������{k�Q�?\��Uqs����".Pbóq����꽴xWK��0�p��JL�.㝰ט,�H:]UEę�Y��)�Hɿv�R��.��A�l�m��ٶ�&dn��#l��vy�u(a�}ٌQ)IN]A��U� |mQ@���.fy�V�ď�ī�h�l���� eò�����=�dB�K�Ԍ�����$���܋��ԝ,���(ޛ�v���0>�r�$��AM�q͉�z̉��G�Jv�q33LaC �$��υ��� OT}����]?��O9�O����7=�(���{��}k<��/�����ͷ�����L�iێ�O�����釁����wK��9�Yt������Un"����ZHٌD��88"b�,	x^|�T�^��b.�``d�V����3&~��ۄG�o0SE��y;Kt���p3�1��Ґ���vG�e��0C�ߴ�͈����V'�g�T&1���<�b��䥫�Y&�V��G∯崆.x*g ;kƁ��J��~ږ��D)z�6jnA���y�����M��J����
5t��\�t5��?Ce���&Fpʆ�\����A���KȠ�od1����Qx@Z�i��m��Dtm�:���0�� ��.�Aܪo1�$ꂵH��}���"!���8cI/'h�n���2����^����jg'CL�uNӃ�����Oqhl�����7ό[O3g���ݮu?HC}[k⫺|���$�[�+}S�У7Ln��y�����-�� e��!���M�$�ѕ8�i޲e�GB@��;Im�?f�a��b���Cvѝ��P��I�i��|�ד���L�	�^ �4�IP6� �4%3��b���,�P<9�_XCJ(��z�Sa��Hx?&��T^����ũ�����mMy��p�F"���v#R�[���c��$`��-@�'ߤ��"���zo�������;hf�5�m��F	�ْ8��IB�MU���e��E�\����%�ȴVɘ�X?�z��H�K!�W&
�c��m�\��=���V�iP�Fn��lVzW�tUO&�k?{�a[��ĔE.�]�R��d?j�	=~�t��뱺&�L��n���9G�|������X���'Jb&����}�"I�G6��@�{ j&F�S0���,������.��j����gʪHO�@L��K+f��)���~�������n)�N.��"�ď�7q�J�(�	E�_z�&z�	9/��|�Ca��>��� @�j���͆r%"%�-:>�ŏ0z0��"c���������T�vt�4���t`\��i9
��@�2�^[�TUGEt�n�e
�3=�h��4�F�J�����1�J��&����*�8
�b{���8V��"�{[Iy��12J�P�wG��c/q�õ4����&���l����Q�A�7���5���
�:n���y\F��)������ɼ4��Bj�kLF�[o��T1'�	�RyK3���U�7��X��q�W����A��2�3�wqxS�^����U�c7�=��-қ?.(��eA+:����hf,T⡈�!���i�֡qA�uɿ���F���nJ:�9�C/�m�L�$�v
}�*�qS�]�v�q�v��&e��c��_�ߡJl����0ώ�b�o��Zei�T����F7J�s)�d�+��劏�������Q�h��7��n���l�����15Pa�`���y�s��V��C����2��|AT�vO�O����0.�G�u�z�7	FSI�eLltbł�_x����)o�U���v��Ӓ��t��LO���Rd�o��o�� $�B��Tz�}�o���O�֗�i[����e������Gs��\R��	� ��/�g���35�*c�ޞ����)������#(���c�@��Y�R������}�_ ��Nr�!	e��K�8s��F=&���sƔwr�z>����;�������XxNi���-��f!�E���hj"]?^��1�7<	՛�@7�.��ûHd�{H�ӊV����>2�'d�b����@�)o�b���=ƺ��su�'����N���ta��I�/N�_6��:��a�h�<7��8��@
���������ek��^~�6��Rt+���R��k$x�g�N'� G!��s] ��8�w����$�9>L������|7�9�zD��1��}��s~W2 0�Wa�QکF?�U��� ���OK��%{Q�m��A�Ϫ�|-2 OK�<�;fOL�b.��+�:���;	���l�6��M� r�;�M�3�ɢ6$��/�E8�#��o��c�[��M��(>�"ߘl�nUXY
��5�ɝ������FTS��a��B��f�c?!�)��9*��o���ta K��U�$��]�"�W���E^��tl���X�����HX&ۡ�(�[�6�l6ԩ>��FN��~Y9��I� ז�$X���v�<��"�~�ý'�0N|�_�a\�����UE��*��<h����7�/�^��ݩIM74'�I,g��Y�`���Y��o��G��TX6�ྶRsXA�^�F��~u���z�NE$f1�B�4Y�K�b�	
Y�������V���q1�7$���+�x$ ���L� ���@ٍ�����B]~t�ǘ3�b�������0�4���e�z_r�D�_��liy�b��^�z8wյ�N0͜$��kù$mr\�݅����,��c�4|�>�<N�׽J���b�����OV��!�<��P�J�k��(��t�ZtS}�^T��7>�pI�ma�&���VɚeXY���|N+`I<��]a�!=���E���P��.\F�5�ZK��I
�p�8W�ΐ��4��C=�{������!�ā��A�
v�%�{�V1`X��M�v$�]�YD�o���*�����!z����8}fᑓ���z>̕�QqG�Q�;_�h��]x����Sy5���@�?)�W9u��/�q	��p�s��6�*^X�D8���]06�Rд��?{�[����hh5�9�4a 
�G�@�C)(Gg��m2 ֻ����0�7~`r�'r��ו��7I��Ņ�ɢ�V���ҧ�{��X�[8G�.�㲃�$��hmk���Q/�� �˕ժ!;��|�}�s�sG��\��T�m��rj�νKT�22�{�L�Rk���+<��rǿ��f^���J�p��c������(����RvV>�mt�������I�s�S�(O��뱫@a���l+��V��
^=����{�+s����op���V�?�.qhu�X��]��ٮ�����9 g6�o�'���V�"�f��	��b����h�^����n��P��>�S�̦��_\��+{}�Cz�����]U��鰧Su����s�rd��f�!io̢��J���9��=�14�,(��-o��gq�d�����wй�f!P���P��.��sb�c<�O�1J����9�H/!�.�{��8LHS��D��T,@�)��!��=�4kE2bD�T��]�͂;��|;���6�BA����E9�w�%��Uo��!��+ZȬ��Y=��,��i^�α �9�$n武�2t�ʊQ�qW=��~�d����+},����{lE�3��E��*B�CI�h��r��-{�b��PPHf����\:�	{����EJ�9���b�� ~�v��.�(�\�+��?���5�B���ˆ� ��˩�p��3�7��vK�����ֵ�(��ڟ����V+%���m�d�\m�43�P1�Aq����_]��}�7�Ҧ���=u&8�t�ԯi�Jw�՞qz�4G�Ò��b=w��rKLG?���K�`GPxS#�y�/Gz��1� ����+0i�l���ѡqB��Ѧ�0R4�������Nj��&�ϟ�Xo:J����ǫ�Q��T�/2���C����;�t���B�#������ť��U���Vh�C��(ϙkQY�j0/xr��O�� Xkt����fТ�x�&�n���,R�+��B��2D�)�ۆ=$+4[q� 8�?�`��?��=&K��`ZD�w�^{1� �nR�n���A�q�7��.��xo�9b�@߁�UA�q�yf�Iα1�h��p��Ǒ�1́�bC�bD��t��Գ��Ke��r���=q��*Im/����x��D��:����r�''="�t��p�`b;\�v�y�$�u�R%�H���$���=�Vx���rM�S��!m$�C�&570L���tzb&�.�%���_���k�E��C�e,ɺ�? ��t�_8C��Zd6RL
C09.�d�[g�)d+H�fj'|��1��=����pb�. ���T1�չi ��p���9��o6�����7�Nd��4������ިl�E��̛�N5p��e&�	a���kĒ��kQ^��`�G�����4�`)������g��y.�U�vPp�nVU���<����a��0: FQv���:����/*�����|�.5�57��� �Q5�g��3M"����+ba�5f���	BX]С���:B�b�a�&��g���$��F%~B�*ڔ�ɹ)?g,B��Ɍ5t�V)��-�Z� ����E�-7-������o�_�sQ��g���Թ�����i�Q`�����B
+$�r0Z(�]^����ꏪF�߆<d9�?��E�PG��/^���<~���ʦߡ���g4DJ�'�'����1
�+�y�^��ȧx��0��K�{DE_����g�qe�<��(ܤP��\X��_�r"�����h��=ږ��^q��N���<2$���������)o�Y1�����D�Œ?3���NN,<G&;Я��t$2��I ��L�ݢ����ܞ@�)bv`���r�6��=�� -"GI9Y�CC��+/��x�$	?��{�e������0O��ܵ5[p�_C�.�yB��vK��3����sHC�B~��I��ux��Df}��������=Po�*L��谀5���7q�Q;��.��a�sq,�	�钟׉�pXLQN�^�/�!r�I�{�W[ru��x��F��*r%|j���uk=O�yfZ��^k�x��	���χ6�l���OY�I��*;�C����Q#���6��↩"�r�2<\��[nq�ׁ���C@��'�&ϕGAJhR��iJ�������5'	��M�%�K�|��$辉��T�$��E75��!��[��[G��4�h~L2�YK� skxm�gP.WȌ����Ͳ� U��ccE}�����c3��R�܂x]�a�t:�/�_���Ϗ��B�=!y������������a��5.0�7_�I����>��iE̡lY]�e��[�e$&�-;�&(��Cmi�8���
p�����?uy�-����-�����:䅏�Z$ߍu�׾)�=mB��Sw�M˸s���,8I�p�6�<�p6���hm	�`�H���<�H>V�04<���7�5��Z0XuR<�
㲧�^�%�\���u��wŶ���L&��<萻� �������j0�Ģ`���������O���?���~ZH�i9��,��*yِ��	C�j���#�>`HUd�#����)�r���8��F�;V����1<g�[�x��!�2���n�Bጠ����U�d�\y���xu�*����gk�N�`�3��DlP�� f��Z�o]J�<!m��Dː�w��{Z ���=��h�<�}��-��5�m�KN�.���x,�uj���B}�0pi3��;���4���Y_�Jz���{d{
;�� .󼯠�F��3S7u* �:B:�-[�u��X��@�i��̨]Ch���2����^
��pԢ�<opl��r�s"lP#xv����;q-���*���ˣ���2�h�]��T:�2��~H��v��F��Bq'8��(;�jcx�U:��?��e�`��rbA6{#�Y��z�>BC�QЁ �9��j���J�<��}�DNڒ=�T������b�ߑ~O��Ns�c�x,B]�}��"�v.e<FU�E����%Y�u�����oSKx�d�+�|�KM;Ch$��Q�"�?I��>�}^uVΧ<��P%H{Jbծ�`����� _�,�m�T[�m�K�]:қ��W+k�5*�
s�gj~tB>E���'�^��f	��C<��]�&���:�L�J.<`��'�4:A�/�k����Lo���
!�7�&�u��N�I4�!!�`���@� U6@��T8�bϲB
WId��i�.�p��+����;�M3����ލy�4�)z$��;�G�����E�.��X�g���U��ϼn�Ȓ}sA�Qs�E�H�p�Yc@�=�_����#�0zѽ�K�y�=�O `�g"�=>�F 7箧�}<�-��̈˸m�y׏�J�kP���U̠��_淪j��(A��8Q�͌��(���p�*[S,-�� 6<�O"¼HIl=�Ӕ�,+�_H{�Cp�r�R�,w�WI�}M����֥��#Nei��?|��wfX̄�/�ۜ�g� �8�d����BT=0�J�4
$}�	8#ƚ`l�j��Ha�eIQ�f䅑�|�L���w}~����n�e�G�^I���9KDD��KaI�;����/�L�kr�=I+jB���W���R<�=����؂�vrB+9�!���|�ۡK�𸟮�n���+��;�ġ?��ܹ�)��>&�4Y�ӣx�'f7�9���篿���!��=�Z�8����0MZ2%�;�h��~�L�S~��x�^s�������q�q���;�7�d���?O�ew��|���&���PH|B �.ᡩ�B�^�r�e�]��q`�X�rcfC�wZ�=�B�OU3\pI;�>2��Y�&�X!�y~�7�S�B �)RM^����i{��	�¦�9^~�#�M��D�B�<��|ԮS��x�!���&��]ɚ`�Ma��g�eS�>"XbVV ������p{�ϦГTW7���3�l��(Tf�O���N&f�E��~ݨJޔOܺ%ϭkßk���q�j;k��qӴ��L�{��0�����p䖳D��NY�_��(�u�[����Y+�5�@�p��w�7fP�>�?1��dU�>�o�d�j��~z��R߻Ȍ�����1��IÛ.��w$������XΗzR��}Ƣ>rA��C"��}+=yɃ��ѵ���.d��F���V`�:2Jː�����Y�>���i��"��ybO�D��^�쯔QLl�%�v�+�pԵ�l~;���<O���+��`�՗͆V��KC����n��lҁh�W��[}t��Q	�RB�g��c�;r�
�K\�<�ԛ�e|��\x]���]Pv�ћ*�?�}������@]��=o��~x�G��y�3���e-����$��v.�ҎY7Q�J1'}�y�����\���ƍn���~�z�昱���G���rd��G�se�Ũ���~���p�A ����k�7]bJ�2���}q̄[�����x0�_�iF\u-�-��p��n} ��Ӄ�����K�'�/y�(�B�»sȱ�j8�Đ���_����<r�Ht��m�5?h�N'<�Ie������� hM�۹I�>�]��x��ZwÈ�����Sh���A����v����xԐ`���W�,}]��?ï7��w�=��ܵ�3���́ omoӚ�cdZ����=���[� H8nǧ�a��;�Z��'�Z�����#o��I�6����U�=x�0f���'�>�����ÿ�Q�0�H�C=�?��xRV;���z0Cp�6�6��*�7p��I�N0EB&V����p��s��<kD7��(�RӗyW��-W�}��������ǲ>-���ٺT��4�ŧpD\�r��X�\����[O7�~)��;T���^y]D�c�K�pQj"|#�m�y���N|P\Ԝ������зM�i55�<K(�%��Lح[�����w��
J��o����ãw���I#�����d��(�T��)8��+D���dS�jO�`v����j '@���}bZ���0ݸ����F�'�cK���JY�f�	���͟�ୀ��]S���ޒӓ�]�
�i��5���i��Ѧ�R�{SV{ƞ\��USM�op���x$�m_U|��B����ޛ	�1�<4��^�(�\��U�<�K}�r�`����p�{�ʗ�1}z.򠍓�.A����M���˸�m{�v5@?"��E�:�m��>]X���������>3�p�����$�j��*�1���#�$V���w5~"�>3��ɶ;��~�-6�~�gX�/�[����閛�}���!��}e`b޾���4\��&�F<k�ﯙW�!�:d��d�[��R��Gk�X��ɘ, �}?��7u]�K����#Y�e�kkf/Dt+W���+
���qn��D���l��:��Y1jJ!����:�6�U�&��G��]�!�4��z�����(U����[�YP��ȥ�ڒ�w��/���I&~`�C��X��������7�F"�_�b���nfܩ1 5�[��jI^*�P`��8
g7�-���:c��u��OL3njaW�
V�]Y��?���\��0������m.�_*I���׼J��m�u���7�=9�PO1h+�ʅ��~�qM���Mz�����Â�+��������Q���?
�U^L��q1�r�P>�d@�`P�xMW��$![�4Tċ4��#0Ҁ��5D/JӪ�O(~���
6�효�xH��27$�j�:Y#�\a�ޜ[g����>_h���;�`�;O��I���z���$H��C�ڡ�h�M���U�&/��ר��9ϐ��!<�yb]+�0�JQ�Y�I%ﯕ�D�!p���W�5δ4���.t�g8��:�cԗ���u��rښ75%!��ϐq�;�|�C��l���k�E C�2�a֭
:���QF�F%_�uQ>�W�����7G:>��|�!/K�v/Jo��5�o��(�V������4������9��q�0�&���c�:��Ye/(���7����@n����]Aj�f�G��~"����8��4�����|���*� �sH�d��������I8�h4R�����3a�
�H���K�Ǭ_��jSZ<,� [�`��z�فZwW��_����<��$P𷗸�R	�C�|���kt%)�k�ֈ.�͛%� 4\X�@yH�!&=$cv���,�B�M��v�P!�[ ��,-t�9�6��>�>HcB�*5<��B�F��7]2l%�7��f�����=kV�Զ��;��juȶ�����G�%4,⼿8�wj�q�#�@�y���*s/[��z7�3d��R^��ڳ��7�"��y4
��š�Q� �w����d�<���+��!e��&�Q�^����P�� �M��?۴��������3P% e�����Nz���8��S.��vj$�M�l,�߷0����5�h��H,�[7��'q�=��0�4�+�vS&]��A"*�Ulv[,�c�|�02594�7���N��1UN^��0��,ٺ�'@��4m��a7�"��{������	��P�OZJ��1�����t����[��G
f���2I�_t��� �v=�����~rw3�TR�dhLXQw[�����*��&ֻr��Ê���D�����ؾw`�OK�2��lI�%2Z��T�Պ`���S��K�H���Ϟ�*�w6�An��3W�>�P�
�b���?��hc��~A��G��U����'-t8��,�Mz��<t�U�����	�o�����HN^�Le���؀]�؆�Cw�?̃��l�T�`��g�/u���h;D�I�5l$��Bd��Eh�8�Ư�}c�c��o\=�r7�D7CZ��\2�!C�"`���_�a �_��V'qywtO�=�V��X���l�B�-B������%���49?�i�q���a>�������?�P��3�Lf�o�Hĥ����Y�'�<���̩=
�͂^����Z0z	Ω�t=�h���ӡ�� ɝ��!�a�>O��gx�%�?i4m�B9�ؑӟ�F�ކRE`^PG�vkn�#�ϣlpO[.{_�%i�8/CF�c@�ճ&t��Gd��������{�N�c.X(i�*bPas��6Ƃ��鶍:	�5T<U������b}V����������/��e��2틻�. ��TÖ3?�݋j��x�#:�mmψ�]�����^��;���'��Y8�%���_��;�hԩ5~:�d��A���I�RH !�[�Q�xP��͜� M�W6��~�FFu��.Ү4���# ��ܑ��d���9�`T���a���'H{=%���QW�iK�-�9`
oW%��$
V�䦊s�8b�@ù*!�;�����ͯ੼�v�w{(�j��8�>XI�O�k�ܥy���|�̚�Y�i*�t,���mu |�Rܡ�A�_���y��vN�T���i���pd&���x�i�#=r���2����E��?=�c�u`jfF����L(\~���1�FJ�ӕ<t�.L+L��^��ڃ0��p+�T����̆�� k��J�_^ƟK�a}B���Ӝʋ�s�/�K)Bg<Y��_*\����� {e�)jע�����������	 ب�Σ����㢼Mf�ߡ6L��D.�̼�QZ��ɹf�1����.�6v��K^�Pd���!dэ~�V(��aR��q)������ml��ך�y;=YS�3���s_�(ci�R�;�����AD�7Ĵ'�*r��b.�C�3P�8��^�벛��	��u,�k�͎�_ ��N�xB�.#��@1;�<1N��I��ţw�T���ܱb����?�R`��pr�V�����	�?7�_d�(|�bu�O�E�b���t�9�iʧ����8���.\���J�	��h,��2&�!f|#�M��~�_�.�-�94E��Ӭ_;�"ѭ�u ��[�J1�p�Ԓʣ�}�Ʉ�TZ�<�?�B�\��0`��Qy��9/d������/��-����/�V���U���"櫑UиU�n�������y�p�'2h�Y,F�	�?ݴ_7=J�RA)9.f���?탮7�����tKN���p��Q[{)\�E*,-��C�`=60��4�
{��/*O��5���R�Mzn\*���	M�����,�}g[�ȇ��)��lʗ�A�h�;j
7��p�r ��c�%�n��*2����h�U�P$s6�UuEU<@��YN=���ǌ�0�*鈺��w�a�f�Q�!.N���U~�
��%�V�������E�Ɋ���w7D]Onk[�X�F���2�p�Z~���O}}�'����@�_��j���P�cRvV�$�
6y����ZA��wa0�V,��Y�֪�t�X���}��<]uF���v��n��C��rb�!�(Ǟ�jy��Sjn����So3)�_R�����������9�q�L. %æJ�}��;���?�a�\9�]�Q'[�Is���Iv���Fx[��QϨ�0�!��҆�3�H����?F3r�Z�W�x�i�tp��eF5����I$���;��z��?�haj�_�3�Ym�H���_��Y�"!^ʊ5���S=�A�.8
���!"QGJ�pW�fTW9[���/S���
F�M!PE�Q=׹��F��*(�NU��D��.h����!<�"}�K��-��o����l��ݍy("a��� }�e�K����-R� ���7�A��o�OHB��,�*��[��umLqC��k%� =0�w=E��A�绩Y��K�*E����O�g=���-h}�t�2b��h�� #fE��x���l��SSk�mX��2ؒ}���TȠ��G�x@�k����A�Vf�/����q�&�x⎊c�����	%k^2~����ure� �����Ǖ��ɉ�.u�z�1mI���x���ʨs+$/ޏi��m:ĳ�*A�7V'����\�1M:ч�$��(�B C�0p�Y\Єt���c{�A�K���R1�p�,����x[RN�8����j9��\��������(��x|��Ě#��ܗ>�Y갾e��kH`��@� �@�Zbu���憣�q)~ʉ���A����"����ﲡM���T��7���%�	�)�(�X��H��y��e�������1̪؂w]D}�x�<��*��v��S��y� �����o���p�4�z��D3�1ᱩ���$��\�Sj�#ƈY�W���?e���51�^�)�?���6l�\|�EP�Qw5�"s��}��W"��X�Zw�^�.2���L���2�=9-�'1�y��7,q��z�х/�Y&O�F��3b�a����2����j���Z��g�#at.�R�|WA8<�+҄)�X��g�)b\�.1%u�j��KS��NR�i
`���[��)�^/s���b
^�^ǿG���.{�h�ԑ��]r)�X����;'�vZ�*i���VN_M9rҞ���J�鍴� Ohf�LY>j��d���2����6�����2�K��t��.�'�����j|�5�~\;�d�Ϻ��0M��%T�#��m�v�ou��P�&�qUS���?�l�|�	1�.�*7�0���p���5	+m�%��m#;}!�C���m�+�F�S)�q*ouz�:�5<l<�L�c�@ ��A��ߊ����҂���N3����8�615V|@�����%�-Au;�&s��U`��tEχ:UL�����Sa���㩳�:+�4hR�S�����"wT��Tz@P��D~����W:h��'[d�:��ZnV+;���Q5�x\�_�0���B*�<�%�
�,��R�br*��I�S`T��mm��
�9N>�!���e��}���Ɓ�d VQy�x�o��qr�*6ޯ��E�}�t%��%���i���q�!@D!o>����˩��)�E�(Ɖ���r�9��*30N� ,'$��ئ����x8�g�E~�N#�ؕ��S����i�=�L���T]�Q �l�<B�_vS"����+G���^�0��{�g*F�����;�LO���bCV)����sE
9�o������f��g��ɡ{���nߙ�r�.	ՠp#ʡ�ϥ뭹�e- �Lǡ�����`���H��,:|��Z����V�B^7p�NH�b��v�����V��l�^b�m(v�\���$����U	�/�$� ��[3S�����'�]ެ�����Ex��Y��?���GQ[��s��'~
�5\�_���l�+�)7̪,���_�K��Qg�쌽G}뾲 #������+S�]xe����7�����Ё?(�zӵ����Gc$�:lu��s	�'tW�QO����c��#zO�ӲP���t(�g?�u�^ojڎ���=ݡ(�����gP�+t(��]��>jn|U�m���%۰_zX!�ո�5;O{M1�t\�1H��a_r�c&�]	�G���u�	�,�-U}���	��I��� m} .!a0ˀ>���T�=J]��q�;}�@�]�}�%�m�/=����TV��F�;�*ɝ*��[�3I�F�B�}O%�]��q��tT���"fC�Ĥ{���d���C�'�:UE������jj]nb��K�WC�t}�/K$P:�0;�]���o��y`r��D�sq��$��jE�TW��b�;V4��p=�2����G8��b�`�|��g^<}��������e�D�u�EZ�TX����~>���.H��V��"��F���[<�����Q�ɡ�k ��k]����3��[9p�.�L��-��l�!���iP��S$Q�D�-(�GK{b:҉_*ހ\��ݍK�c�sR��n��kv"gC�~X#Y�c���9Fߴhv�
;�mskљ8l��d%�|䈘]�6T�s9�v����VM����;O�]v�;-����U�Gb�u���
'�N��Oo�wjȞ�����[�)U��!��ދ�w_�Ш pVB�Ư�*>4�D���y|�n��)@�Lg�좬��B,͇����v[��F��	Rv3���'�����?8��ُ�e�*h�뱋"BY�_�fFga�؆��z��RGBA��W�^Z����ƃᶛ�7o�<�Y�m4��\���U�����AZ��FG��M#	�VB�ϔ�#�$�ɘQ�Z����9�>'��$X�;2�I�Y�}2��K.AIk���)67誐;h�Pĭ��m��-���K�n3<����.Lj	0��OϜ�<8�UjZ��N�f)�XA^��J��ɔ��c���w��^C����Y>'� 
�,�x4��7�V[�nQ�E{��\����Q���̱t��Μ�	Z����Q>����rK/q�5����ss*mX�q1e��hH_�A�&{=��h���-��M�B5=q���Y�SrM&��5>$� }�(6>���؂�"�&u���8/J��Q�q�G��P���WEw\`�,NB4�O/_�I��<����hk�B���r�Yƚ�`�
��p:Օ>�����p�0��ka���y�
%�˷�v(�+b���lFu��jvu��;�t�$�]3O#ui�lu�I�'��Ōf��ϲσUa9�[�TT���J	)��]��a����LT|�7��qxA��H���c�X�/����g�5'�/��ڃ��f��LZpd��ZTˑ�=��o��3�&�������2;�Q�e�#3�mB��ht�'���w��-Bx��"�S>B��-S�F��ՎƯ���9���j�m��ԡ+$SF9�}�ޠ�%{$L��Y�}�-C?J�8C�P�H���P_%�]���C��P8!2��L�ȡ��T����j�%FY�ioN�W�z]ήYmg���)br�/X��60ةV&��]�OB)J
'MJ�Q<I�F�D�<�Uv�`�I��H�|�b������ɣY%VU�4��,�dOئ�Ab:��k��eGZ��2	��*���������}R�E�>l<c��+���C�$�Y���	���ݞ���h�+TT�*֛e,�f0����C����WֲMWxv�z��q_e��SX�-��&`jiԩ����{U�%
~�Q��U�8#ZAR����&f�j�랸�=�Ff�*��If��2|�dwS#�������vF�����r�G{c̵^`w�P5Y7�ԩo��R���8�-��l�֟J~E��U_�j]aǝߩ�$W'}�(R3t�G�ѡ���)�़q^V�Fa��Sԍ��n�2(�8����]�V�k���2�F�͕mLü��Љ���V)�֮y��f��5t`H�Ȃ�E�֯�a��ꭜ�.����6����Z�b��{>�����@!6˾�x���`n�m�JW���2櫃�j��i	W��M5�7	�%\^a4|I�����p&�=r�o���/M���o*��E��+��7q`�jHLNw�)З�����icL�4]m���P+��sx�V�U���A��b�ɝ��A�z�p�����!� ѫrx�%�S��_������Eݤ��Jp?%ru��i$??�˴� � I��&T&a7��
*��J��k{�C��[2L�$w�2��캇�w�Rv���x%�R"(jFf�p>)�s��⊖���@,�=�U����@@u�8N���d:!��c/�	s�}�J�*���Y��\�B�1b�xD���m�sk�O�5J}������%:���íڟ�J��m�(~�kA�����t.V�Up��ʢ�E�e��yX�r���SR�=�ʛ��N�%�ڒ��8���QWR]��Q�T9켭�!���f¬ �[�˙�lI�@ �2z����\f�����4��-�M��D�p�B߭��\�:S'Wr��a��t�ϐ��b���A�|�s�֛W&��ص0�"�B>Je7|�hpN*�\Y�(�����wb'Ų�9L��<3�Y����]���Ğ�B�U�p��S�(Z�:A����];���A�[��~t�����W�	����A-����[�@�����]3�V�J�kM��Pr"r*Ag^���Tp� |��J�3�E�n�<U�&��}r�t'�D�/�y��+��-��"�c��@���h�L3������&X��=w])�5�ή�`m$,l�.��q&ϫ�R�z`�o���� h���v��,"�vy�	�zc�$:!��j@�}ȩ�O���,�R#�2���yB�cf�2��qN���0ZR�5��B���7�7w0e:���v�����Ъ]�L����T�G���=�tji�����>qC��B��|n5PM*J�dL�˩%�twU���;w�x��6�P;F�M���B�Za=�4�A����ٔ�1^�Y��!�x;ڟlk��(�9���)?��?W\�6��&�8��؅��R��k�����$���;��!"}Hh��.gٜ�44u ��&5�:9͙ǼC7jP���0tD��&��$8�DO�6�^LT�J�i�r JN��oʗ�0"�9k�/��iC<�i��;s���<��~�F�X�Kp��C4	εɳ�/��>�Q`��uēŜ���[oF�gr�\.C���_�T"����'�����%<�-4�q�
����?MiÈ�<�OF��{����Kw�m���]_iW��cj�p+��
��|`�5�f<7���7F�t����(��G���*�n�n�gz�Q�Q��������>;E1�*�?i|���b����a-��ͣ�h���8T�um��r�jV���|am���<��~��������H��vb�����1�Äކ��U �-���57\N`� \[�9- ��G�F��;�5b��L>��{�u����e� �J����i��(��_4��~�����a-�C8!��A�s�>`�b_U ƴA����w�V8��&ث��#�mo��=��Ҭ���Q!`�C���Y��,A����E�ē�t��&w����M�V��qp�8�]U(�x�>4ҘBǚ���~j�h�Xt�_~��coW���n-"^�< ��&������	����׷��KS$^��<����Kv���"�磘��A�2L���s��
��ua�}[��"x-���A���� �7<Yt9���H �,E�RQ{�r�D�cf��a$���v��6Rڤ� �:uI8�8:��qܔ?�ר�4��6~���jd��<?�;���^�����(������[�hE��F�¤�3@t����Pv���RO�RtD��������M�����T�	�Ä����K͔��ZQ��0�7�m�s5�aR�&��Xѫ�ϡ�	�.L��N�&��=�)6W��ͤ��B��|OB׀z|"А�d������e<*�l�M��?�~�x�#����xe����Ϙ��(�O��s���c`����"�P�GsI�Z+��5�4��k4�[��Y�7*��\�{\;��o�V�ŗ����W9���k�^�`�4:*^8[F�T5L��/��H���C��Ba�iڰ����'�Ŀ𒥞���I����E�U�j5�!v�Y%�i�~YJ.��2	�SPD�˃�k�,Ly7������J*��Nkm�ٙ
@�قl��=�����eW���'sUHC��n]Q�QnVG��j��B]�6���5ɉ��_�0��ɮ�����&q-6��������s�(�\�OvuH|͕\U������3�TT,�O~���䎮?t��.ZOu>��˕h?���Uc��y��{�m����4�c�館���c�v�:'7���J��--yg��Li��;�G)$�`5X�;���\�W�H}�譬�y�))
Fq�N�Z+�0�h��{���
�+��B��[g�P:\M�Je���;?͉'ɅYjJA"Ȱ?a�f���������K���t>��.�;[��+x�a�J^I⑻{�v�Q�2
[�ƿ\���r��d^Rjg����7����b��B�Ė?�9������Y3������. Jpݗ���#�Q%3�}��A��4g*��'6�%�kluV�+�7�#Uiv�	J��.��ĢG��^�d��Y{|���`�.�.��S��]�R�~�9�=�A>��&�q���O<��4�oy��v@�Z]�������˄��JeΌ(B�F�GMtJ�6&/�ӂ�i��a�S���3����Rp$�~����Ӂ�֩�	�q�엑�:Ihw�zE��ps�q�s$�ӛ\J��,&�?��>k�����@5���G���+?.�fv5Xr�sa��c�sX�0�.mߗ�Y[~j�%�|M��M��2`e'$�+)�Z�(Y@�����"�r��b��+ ��%X$]������ܨ���Y9>�c�{�m�:���V��=s� �ռ����לLx��!ft�K�,e��00CfbU��/�y?�z�_	�UV�����=B�K�!�W)���X�e��[��ͯzytP�}�y6���y���}����,y�>��U.��~f���{�b���$���k�Z~��k��,�.��])b�d�"������|�_Ԡ�	a7S�U�R��ğ��m}�VsH������Ys��Gв�QJoIl_���"�"6\��C����{�d��O4��L�'�@'���b�
n�s��XZ���p�p����� �:p����H��W�)|y3���λ`gX璉��ݑ$f�@�!��l��WH�':rn�:Uz�u9��0�~%�|��_�,��Q�C͆�<�W(1�����Jm��z�5�`8��8oܑ�!QƬ-W�*s@HG����SZX�)�!�w��oP�l*Euy�pm��\�|N��b�7����5EN��1VDy��p�Q�.�?K��v���z���34�;%~����unt��AЅ~�p�b^��jkg���}�=	d�o�ЈF-�O�����k����̀z��Q�TO	u�2Lҥ�|���jZ�PŅ��-�dg�2���ޠW��6�M�n4B��@x�0n\��S���Y��D��Z��Kn7G<F�;˵�T�5��m�t�v�O�a�Z���&�y���J���2���e�2ye�wf���t��/�>t�;W��w(`"�oh�7@y�b
G�J
j�L�����T�ڊI*���Z�X��*�%ϰX�s��|v��lK;���Y]���;>{hQ���[��ۦ7�]gi�����'u�������{��#�x!�Id*" �����|�%���_�xY>�gO��W�^##�����Q�l7�r?܁���^�--� CL1�&e�nw�[������\l�iBYV�Ӳ$��F���>Q=ea�[�� �]�5��
Rþ.g��{��=ah�5D|�Ʈ$�s�A���1��:���7���ƙQ�]	ҵ���о�7��pl��y�с�W����8�1Ƨ���X2pr�`\�2�R��p��ó�9�+o��W�a�V��P�Pr�
|XA]�;�r��>P�$η�D$����4��G�k�A:�q�[���D��*���J5 z�f��ϛh/�v��!q]%�����۩�}J���i�܄P߯>k�>h=�H�U�[�|�Ț�S��b|�sL$þq�0��X8Cw���S4D�wE)����e5�T�w~�ӛ{T����\�|&w�O~�% Om4pJ'�$���"����uE_?@��B>`�Q��WOg]�;�<�P��mx��g��R�tQ�o/@���(��~bZ���C�A��4|��>50=��/�)�T�"=91@]�u�'�*M��n��vF��i�@#�ݦ�Dڦ�����km}��%��������䘪u�Sz̦���Y<K�,v�@��������|�0dG5.yc3Q�v��Y!׿�2�u*0`��q�%��}�m�BĶ�lSܯ��C�MA)*�w�f�������C��~WͲ�&�A@X)�4 u���Io@^L�a	�W��r�~�\��������!����y��� ���
��ZP*?��F��{!a�r8ň��RB"~�9�E���:фs�3wbbB-=��w�^>��I%��\���F\���w%� �����#Xu�\���LĹ�a�th�ق��{[h�5�9gB�&�Y9lw	�W
���O>��S�\?5�(le��{�9�e��,'��f2}!�*[�lG>���y6�˥�PJ���=Q�OEA��z˹-Vg�qK��t9�FZ�#B���
Ϯ?�c���c�ֹ�8wb`Q�Bÿ������S%l	��ܝ�;��������w�ߘ��j-ނ��~:Y�0?Օ�#.���-C�C��!�z�$���:�_�Z_�r�U��[Yn�އ����Q؆�Ɔce����7�S���@���/9��ϸ��2>�A����}�}�*m\��oV����r��ifۇ��M?R�jRy�'e6
�ܝ
��-a�՞���XNߨ>��U(qj��`�I.}w�B���������b�jF�&�٫爕A���T�o�U֜���@֩͘{u�S�=���=)WX�SXfw���~��E;�w��!\�z�	He\��/X'��#�����^b�z�G
�>>��K�Q:a�O��y����{�=�}%�<�@��DW��B%"�&L�ec�����^)�*��%B�ޡ8iE�}��?Q�S9��N��cAZ��Խ">�cΛ�T�6��o�!����7� ��V�CI�Mm`��kȪ@�Q����5�vz��M��y�s �����
N�ҙ���(�0[>'�AG-������Ug� Dk�an�kcr������h��I�)/�&J3�;ɫܑ��Z��=�#&��!��"�@ͅw���c�i����$�w��j�Z���Ζ*�
��6~��Wh�,^��o�f�ܙH�����4���]�c���|��Q��\5&�����w�SZ޻�@�Lk�k%`dxDc�t��]������� �z뚉bh�/!�P�� xtn]=�ʘ��n�o�]͋��
���-0�hi����v
����m
�z��#)jTtr_g3%�����P3�������k�靵k�x�c�̼��mQr��(��ͣ�~Т�/cV��|��&���e-d���k��df]�*9Xg�
���O�W�s���Dɹ5�b��:]�A�ú�K��;�����!i[�v��8CkӨD^Ji(>�'n3��ѝ���� ��lKJ�
�w}y�&��ԜOĘ>�ӽr-�����q��%:��V�ó�*�L��"c��]mf��9$A/��8X(�$��U]?4�� Z�`7���x
��a���j��8� ��[�]��Ī�Ȋ:�Nt��IA=o��Q56���KXS�8��̈6=7&>m�F�Wd�}k%ݕC$a�/���T�Cc1{!K��	����#��F��Q�����s�_P�
D�J��� T��J�,[C=��e.�Ύ�����{Ǎr�Ħ�;�an3�[���7�,@UMZC"��j��o�U��i�^�PK�e�#��;�Ұ�|��/K�!�Ù�_ڲT�~r8��R-ӹ�I��z<�.D݆����r��ז��O���+kr�2Y��xm�=�"�)3�!s6R�m�I/f�Ҍ�\��8 �N�km��Oo���k�
��@���� >~u���:9(�M�e��_�'x�b�ߚ��9���k@�Ind�K�˷����2k�]+9P�.���"�����g�	$\+�Ub�8k�t|coσ��1���LO/)��B��ट%���^)���-p��#~�0g�	��|��Z�n;�!j�6x��qD�4v���O8��m�@����Y5�zq�'�]p�W;�m�i2�ޠ�3�V$A�	�B_��W۳@~�� ������y�*���� ���T.Щ��۾���{WĻ����SW�����i�U�T���
嗁���-��b�f�sr'&5Ļv�ZY.��}��B�u����.�b��иgJ\��ɬD腸��n��k;�f#ԁ=�g�wl6*ט4�BG�~UZ}f?�֜5f��jZ��,Do�(��y��1�I��n��|��qBT�v+h̕��U�?/p�H�O�bi����+�V�G���q	Q!X�:��/-����?�D�GA X�-�@DC����N0�џ�P�g�U[�n�J.ˍ�t6��g�Cy�����ܻ�](M;ը� ���U^���FzL���j![�g.�5����)���	��8���� �W��I��������OC8e����E�bs�G&J�gVt��Y�� SX~�찰.f�1t5��$�������7*���l���D%Tf�Im�e+���'��S�͜@eB*�Ք��&�c0�!#T��ic�����ǁK"�s!ؼ�վ��E�(���)޵�����\kbH��|�d�B:h��U�;8b��n0�}��s5�a�5P�er�R;�nJ��软�eq)����)�-� �x/���z�P��ހ��AE�a
ºhF���P"R�g���9���R�v�a�J�# Z�k�^y��x�ZN>K�S�KGt�/���@��XX��� ��N�4������N����ӝ�]�O�<?���80!�[K����$`�����U�����]fF�K鶶]�oG��'�
.4z\_�Ãu9�=�9�f�iK�����eN={\K}`g%H���?ܛ�)9�)��ŒM[�b�BO��1�d�	�NQ8\�1�F��w/˫SF�����l\y��4�����M���H�ܾYL�T�̽��&��S���%��G�'�q�r4a�<CMZ2�@��O�.j10�Y,iUf�g��	�z�����m�z�s����e�I���Ȅp�
�&��,,� �m�W�-'~@Vgc1cjm�C��X���w-t0����5�h�\�.<sae�nX������P��6߶2��n�Vkz�v����X�qr��Uu6k~\���F�c8Ș:�F|���!С��A���IvgÃF渠?^�D��}�4���݇B/S����bi�6$�ؐq�j�"5~fY������gB��!�!��e�o@�L�G)g[��G�n$#_
:�s��~����B�j�X��c�E�'��Wջ�؂�z��ZI�*�K�ТUQvO���1��a�:���9�2I��"��Ff'a[7�M���Wl��N�~�2�<J<c�����=��4uTWB*f���庲Wb�M.lT��"�) �)�Ѐ��#w,|hewD(j��L�B�YF�����z���YZ��e8}k�d����m�T1��y�-%m9���[�q)"AS��t�P7[.{)m���}3�ܱ�'����~|��5@�U�q���8P��nz�N�I6;lL�ͽ�=ؙ��;�R!tA�Ӿ���Fcq� �;W���=�%���R�h��4~���}- Sv�4}��#���r�|R�鷊97��$e���Ŗ�JJ���<����[���~?Yp��т�G��-��ك�1����� �7nX"�AS���4�����C"��Bh��G:QG �Y~��Rg��l�2$<�"���B��\���j��^��0,t� �.��d{�[ �8L�k崗=����A���wh�M1�5B�
�u`h�Y*#�����!ؘ�Ɛ��B�N����`0k}��b��A+�qƁ�Ԟ���� vc!,�ދ��-���Q6���|��"RU&��r���y�F��HVw`���&���L_��2ۋn�p������x�����)��6!QcL��Y;0'�{�i�w�������ay'��]�"3�D!�� &Jm�ԧ�G����n��N�V��U�B��*� ���z�̈́]�:@̼;�U��Dċ���
u�٫sD�Φ;0�,K���ǩ�D ��{��I��M(�}>D
�~�|vf�0~>G���r`�����ɀ/1/�@.����/�	z�;�>?Ϗ��`��e0�ޖ�'�z���i�&�l f̈́B�X4me	�pp�]�f�H��� ����}K�����2��j��1:�?\S�Tq ±��@<��a}̊2���������:`�f�����Q��U(PL��:�I����_Ѫ��[�=��[�S#������M��K��7߅����vy�߀�L��x����
�A�W7��O6�ӈ{t4��E��@䔎ۻ7 {��V��3�ېWȝ�,��a?p��Z�'F��Ntl�sbB u{�$�|�q�-��O����7�&ɢf�~F�����)Ԯ�QؙT���e�����R�ģ�Uz !��l��X��9�7h��iUygBA�m�@�:��Q&Q�v���iXH]+�&��:��M��J�����g���i<߷ˆcn��E�
�:�~
��#މ�[����E���A)�2g$7�nC ��icD�Q��x�J��m[��v�)r�U�Zf���ŏv=�'5O����(��U:Ae�0��C[�l��@��b���xJsP�b.��i���A?����A,5B6�t��_
����ᷦ��\���9G�+�����	s���ֹ��,I�k �N����;9.����Ur|�lyd���⊆"��V�γ���@Si.�~�Z�lh�9�v��8�PB@1	�����R9�?�؊^��Q=2��x)$�t�Q�c��o�����N3X0K7>>#qb���FR�&�]X���d�o�<*g�7�ݳl�$%��_�����a�5h����)��Dݫ�U�P4���E��:�t� D�o`>��"}K�sg�B@ʝ>Dc�����eG^ʭ��M��
�/Z�bQ������h�zfft�6�YLs��g.j�ɋ�G�f�p����'�Ma,[�c����t��A��6�+DhP ��E�P#
��A�lb��1�д��_ ���=3jƁ�a)S�4#%L�~�>��)�P,!z��A�"
X<k�����mӟ��"�?ty���2&]ɐ����cz�%����i���f�q��j�~"8i
���Q$)]����Y{�6T�����v~�p��l�Ɖ&�)����1�}L�L{P�blLH����b�7�QT�'�% zi�?ZKSƮ9B��V���
JBq+���8�أ-"������Ԣ��߬����*L�<na��sc�`9�����#p��W-j�cn�Zή����4
i���%;w����k�sϨ����ӓaT-5���������ch��*Y����[�].(�.����{�~QL��o����gw���6΅��=0d�[����+����"@w�l��(���dΞ0��A�]����f����dHb�P�C�φ3�B5	�ظ�߼�ˮ@,K��fWj.F��w��/�� ��~U�{2�]w�6�8��}UK�:�Kx�����v�i��ġ ��:�;�
��@%Ǵ��/�����������0�!Y-����&�>���B�������)�D�Jph7���� A�z�x�@�&J6�v��S�������𰆀���l���`�а��������yF�)Px9�⠃�ж.#n����2؟�tň�EVS��%��7~��,_ը�J���R�=/|�Y�Pl��!jf��?8�1��2ء�g�e�@�6��zӫ.oH�PZ��K|��)�"�E��|_颌��˭��v����X��iy:P�'Vx��\���<n��'Y����hh��n! ��ڄe�Yj����iˮ'�_{!��R2�ͤ�1#q�D�Ff�]m[��	���L�޺r��o�ۑ��3�7P�r��I�BA�i��|�o(aGT��4��f���J�Z�fr��{�*�]׬�N$��>q�;�p��\�t�R�����|��Hک&���c�;Rx��`�45+i��k3H��iʌſ��@q�	~qʑM��4�a��~�p���l�Q(C��O'��ÿ�_��'%t�C.��/Vho�E�F��QoB�E&��|�0�����m��vo��z#BG�|k��E89�����.�ҖV�T)�r��<�a2<�'-s�t����{��{���OLc9dyD�`A��D���	��-*f���n�����ѿ���;\�m�n=+�>�A\�7�4��h���N�fv���+L.�T�A�ұ��p�WHB����yl$��$5 ��(�w��j�k��)T�J�Fhv���]��v4h)��:p��s�@{�[ҁ(%g���i��Ĺ7��lB����֮�Ȍ$�E��?o�ܷ�T�t��My�=¨����o�������:H�)�ّ��Ps ^rػ�c���GDj��[���sK,��b{��?�&��������
_C0}�1�D'�َ������V_�	����Jt�A�Hr����=Dz"���"�@	�ײ%q%D��<�(&ъ}p&������q/�j#��%b���~���a[,����xR���i����VZ>ɳdh��N�^-u^0�7���a�������r�j���� ��.|/�K�3��u�(t0�� �[�*A�����HW�I�_Z綇xa�,~Cy�~:�����c���5�u��T�T}>���z)���7�U�������m'G�f�2a�uzwnx�=�!���`�G��^nE)�]�>R����RCXv�1���)aka�V+If}-�� d0H���}�t����[��-w�~��B� )�s�)����AM�s��������cјͷ��1�Q�$�Uut�_{y�g	-����N�� �(�'0�2��}���X �.PD�RT@Vy��ˌ�m��a� A#,��PD �RҚhxDM	�0�r9SE~+�2+6�SA�%�Fi�.����'HOT ����s'%F��ǀd�Fl/��V��1w.0Q�_;�Fm�t<7� x�lj�7�Nx��}L��f�,R"���ћҮW���R�A��x�.��!�6���=\
�].�n�e�ac��Y�6�Cz�2=G1�c��9�w�*"��<*�[��b���k��#@m���U�������Z�b�����7���m4s교�t�L�U���Y�=[�"�6��T.�Qݘ聚j�N5:�O[�.Klƴ�v��*�����%�;D
�h��%`�I�*�Z��w4��~R����0��rJ���,�4�F���0k�e�[��c|��N��b�B�v�e������f����G7�7������6l����L\���׍G
�[=yL�`:^��,
�Ӹ{ϑ\��q��[";mm./� ��u�\�:$FZ�*Ab���
]��J,çġ��f���8�.��i�T��kQ!2���,��:Q1ft}��r�������4""�3-+u��7�!.���ÏJUo�b.���[[��!�Ue��1w��Az)����|�����$Qӡ{��=��+�d��qM�?�y��*	lR�8O��QM*_�)��ܱ�|z�mC��7��H;������2�R�+�޾������,x=��n$6��.�o���z63Y�O�2���Z|�B��*��$�Q�R�k��t!&'f[�`�[�o�hf�=1�hߝ1��SRsp���h�ԍ;�2�sO~��i�ź�J.� �%0ŵ�[i�\��ePX���|2�� ��Xt����ҿ)�KGS��ڤ
y#�O ʆ#$9mV-���sb����U�G��L�9�5��.��x��_۶V,�=W�D}�K7��mS�yt� �=G����N+<��kC��N�ʿ7s,�~i+1q��j����k�2�>̩��B���!v���ݙ(�h��\{�P��i+��#����,��'g������DX�I������k6�!0>O�	a�:ӓNH�_�Q�O]�4[�δ
<�c���m����&;01����+�!D�3�C��������J�M�nx0���'OK�O�6($ώ�D3ω�@�w2N�$D�b3w��N���I�)ǳ�N��aA��"���k��w�W]~^��VP)»�sD�� C?:9-��NMf���1ϝ�|D�p?��_Ax`�8'���3<ݗ�']LO��SRKxylm����h�˵��|�RB<sJ�"6�r<xq��}(��W��瓱Ն�OE��5��N��'����|�BU��8y�AD��O�R�9���a}�� l���Sf���S1�Cԯ�5_�]�T'L~
)�k2[@����֝��&��o]Ǜ�톃Z��q��h%�0q�/�������	%�o��#n��z9����t{�a~�ԭ�,#�����,�c��U�on5?U��-�?ML�F	�2>tN|д�X�D��b¾s�7G��e�X"�����ڼ3��{������&��ӥT�{��U��E� ���f��oM>W*fp��Dc�<��<��}}_ȁ߿����8�
���l�ӞqB�[x��aR����E��O�n���\n���9��1�Ȝ�y�u�~�Ljvx������
����F�g���M��dB�SY��Ó�EIq2�J�Vc�z���n垱O�5eB�C^���4�V�֤v�(s�!��s��X$y����0J�m�x��}�wm�2>����6�-N����	x�+6�� eI��]3a�������6!�b���K�rLǊ��G2��nr20eQ�v������(���j�b?��v���z��Rtt�x�!�'�Ms��m�����탁���X4�$^�)+�!wp�0�
��7IZ��T�]�q�B�i4���0�-��K�s��g���2����D�9�t���G���z���vTa �1��ڤ��ϴ��4�V��Ԑ���\m�ˠ]����Bᡥ�Iē` ���� �b��8�����d���/�H�4ﾧ�D=Kж �S�����[�ܾE��d:xr�4#|{�08ŝ���0��;�/�8+�%�`MH��ݳ���Ƽ �#�F��V'ڄ#���*6}��7d��S��;�*�����ig����WcQp6�Laf�� �pgs���X��I�F�@<��Y�^u�>�*Tc*Yua���^Gke��gYf�l����
��3�nO�C7�u+R��
�l�ћ(��|�i�ߺ�#;#|�g�X�����xoZ8��8j;L��DoJ���z�և������.���%�	o&��F8��m�0����΄(:\V��ψcj��=!�S6��V��^���֯�a��;�F_�� ��6���֫q�~���K�c�vB��\k�����W��<jB�u��E�������m��yh�8}Q5Hd�: xU0)ӱ��>�_p�zN�F��2��%@�xӺ4��
:w]�u,�䘅��od�����0�-穩b�K�'cE��� B��P��~��u;G��c���r���F�Dg���:��:
��?�����r��v�)0!�tVƸW��rs�P�I�K�.�|����+r�p��Jw��i%-S��u:���Ap��G�
;W�E$~�l����8�=�.]>ⵅ:	5ɀ�}�Si ��᳽��9&���_��$������B ���~�H�p���"j�dy�=��2�6H����JYCW5��4���{L!�� ��Щw�m4���=`ɐ�l)Wx�w0��t�����cf����O�(�:`rG8P"I�B;4��/��
�>"��f���L[D
1#�c#3x���u�n���F�E߭r�W^�]�p���9�*�IK����A�����5�I_��jcb5���B��T���X �
^��k4��Ts�-�o��G�ː�.3)�IG�l��,�HR7Pm�<�u4VF�x�m���a�(�ʵW4ےA���y�`��D��l����^$$"�A������ڳ)���ݴ�{�pYήvuu�f��2�S�E��O��<�G�#���#�A}�'�_�v���˗s�"��<�Y�*��=��C��1a{jQ��5���d�:��Kv�c�C\Ӏ�yP���Z���]�n�B�mR�d2A�J�_��

0qz��R]y]8�3$�e
7��i`	`����X�A*�;W5	�4w6�no!��6gM��<������Q/�G��w˱�1Β���g�sh��o�6�B�)�o+���t�Y8�~�w�1��?_ŻL >�b�IYKd�p��߯�k����#��9O��+����{'xKY������9�a��Nv�&���h)��[ �A)�w>��5L��7�_P"�DQ�M�m�G�LO������Yqo�-zR��AF�s��Xҗ��&�l�s.�y9�rf��`MQ�|���7|��H@0�� ��xH��Zd�t��ę�h �-���Ҷ�m{)��2D*Q�W_�7�o;��5��P;	��E};*� (�`��N���E7���#��ڃ��FZ �wo���\p��p��z�"�#:�+CpY)�ٱ.�Ԃ���B{��D-���
"�~�v���iY_��A�o TG�Ԗ"rNv��"Ny�� ��妈|��ң(,���#��B�L�I�oA��oq�1�y�مAS�0�����B����� ��0�Iucr+#�#S���v�{~@�����vR��c)3��l�a���'N�[%���ǒ��q���!�*ҡ�@ *U��E<~F}~�〽�3���p�����_�o�����]z^c�J�է\U+����@�4����]UBvȽt4q P>��l߮VݏJ�$�׉_����p�c�ne��P�iA2�g���T���;v� �������v%A+D���k���� ���F���f�(�eoP\�,������t�쬥�R ���V�`�Q�<"3����~�1�>V�4�W5:����%c��2z8]���t���/����O�11����v�dUP�Eف@�J5��>p��ܥkU��lm�L�7/�`��$�P�"���`������j��0˔��Lq��ݝ�ԛ���3��<�J;�����&��_�D�G�*=I����t�o�"�GK��o��w�¶���\�F�ص8K��!�O�ͼfX6�������v�>�n��De)�,�r�J�FԈ�Y�����q���4g@<�p�VCh���1؁�@���y�~05��� ��<�O�{,F:4n�,�<�{��Ty��7n3�)n��(g��a��QI����(��u*���밤	�d��eqgu~s��ķ�^�^"�!��e�9��/��@04*�D���2���e�|��`�ߢ�$� ������O�d�pb��'��>���3��'��3 ~<z��	�7�.���H<vk��EK��n6e�^�g��ó,엋e�XM���)�����tОZʶ�Qj�����	`�!(]Nԡ̠|�� �vC,���霵��prEx 2E3�d7x�$�w_Ѷ�s ��`JB~��K����)P����o��~ŉ�]��6°��C=�����4J�aj�A8յEgܽ0��F���Q9ˈ��]�0J�ax{�;��M�k�TR`?D��V脏�!0]����m"���7n(-H ?.�2�mU㕗��x�};�)�!ɞ��i�� �-4�\��V��ߊ �_�r��+�n�:��Z��7˃��UZ�A�a�ӜQ/=�6Ǡ�n�u�5���Lu� WIv8���P
;�˽�r�ᘸ�й�.�x�K%C�z6����eb���_�顇�4�yv8z��΅���O�PWC��q��j�H.����-�ltO�@�/��>h��k������nuvG����`FnP�&�[O1�9�d;>����>79�T��xn	���X��W�zXD�.1��~��r�g���#��H��K:�Y��ы��O&�aqw�7R)�<�W�t7����4�|�Q�gٚ�f��o��u�0��<FD'���@<��^D�<�����*|���u��:Ue��1,0�Q[�R,��7Od���$�/��EaIį�ƣq��N�+�X)��V�6�\�;���Y�qt��J@N��}9���͝u����th2��O��x�;�w� Bǈ��&ZZp��A�xf�����7F�H��Ȣ �={8�� ���o9>����ԏG{���hlfH!�Ϯfr��#��e�eE2]@��^�����&���]���Oܸ�p*��9þ�IX��V ���I�$��Kˉ|B�ɮ[�[^�S��W�w��;�������`����|��g<v�7�̙�r�\<�j\_t9��	8���ވ"�rj��}4��+��_��^�w�p����Gc��5�U���̍ML��m���Dbz�Dh}i!,�/�eg�
L��$4�p(�%ː���`��)F�����׋0d�ޅ��0�T����ҲT�#��Ba�?� M�
��L
%�='DM��)�XO�5M-���Μט��!��U3�v+�ce��,�7�Z��3�FF��EeM��Q�&�}71��H�ݷox�N޹�<�)h���xF)k� ����^�͹��بj*,�{�/�	^��(]��T�4ۚ(��P[�h�FXW��
�}���y\'_�L%$٫��� �ȷ�x���$=�W
�],UW��2��ܞ��g��K�֊�b�..#z��X��ެx�%z,>��
І݋�7x�ҿ�>f��?�`�y|��Ec�e&Ī��N�*�P`:<%�����_iB���o�,�u��H^��
U�;�]�m���w����z+�^ �I?�)����W+F�a�K��������P|Gel����°���z���ȥ��>���_����MjN-�~��gZ�t�����ɡ�3��3A*��$�0�o��p2�ߩ��1v_.�m̊Nr7���-�с�<��t�&�d��=t4���d����g=��#�"4��S�e��]?� 7�
.[ڹ�����Q�o,�����	��������t��D��l����q�'5����ϑ�r�z�4�8�˘GH뱗V��s�3F�Ls����&����4}���S�Ug�Vf�����+�{T�P��sm�V�Q`���\ج�J����M�'���V��U��M�e�^�M��]9aHU_��\�.��8.�^ʪ�Sن�<�}��x=��*"��ǖ����ɟU4;.����}Zh�_�wXD1���x*���a��=Ds�)og]b���Y�Nl��"��f8y҇s��ws��[�ۿ`x�ꑭ2�����iD*���~q	�b�K����|����p��,2����?��=F��&�l��;�dFv�j.��s���{x_��	ݱ
wbb����"G�\T�/I�\I�J�}"�8X+4��1��D8�G��v�F��6��]K(��
���\^b7zkz�s|��Y�IS�d�C�W�^A��x4�_!��h��:ag� �M� ��a����.ϊQQ�y5�#��@���`���-*�׭��.���>�aQ�x��p.�U��%ү�^�f�zn�����\z/��� ��Q�(�=xm����������w"	�����l�����*��1�ϕ�Bȩa5Hsyb,�jB�,d�5xv4)�U��k���y	�va)�lc��L��'��(=��hB
07��,$$������4�Y̆�gJ�d���ʢ��c���_b��g|�O��V;TnK	E��/��n��]5�\�lS��fB��-�b,G)�r�y��y��R��O�Xn��,�;�������SƟ�	+�}���A$������	�\�׫{��il���$��c�� �G��C���PY��U���Y�I���B�i�^?�a�j.Bʡ��,��M!�y�'���c�%N�`�6s�ժ�מ�" 	����M��];�j(���B��cU?ְE.U�[�T~���M�q"�?��;�������M���cj?��o���_+��-��{Re�Eŏep�P=|@�+ۇ�>��(��^#�ӷv,J�r	�����f*��'Y!�\�l���c[���G� �j����P}㗤&t��- וr�mPd���?�V�vQ�,�`�b��;(�����`����%�y;�n�hE�U�P;�|��I�G4ȷE˙
bm�ì%߅FKO�/�?[ͺ�4��>�O�:���<L^��/�/��'5�S�}�+PUzpu�V���WS�	�9Z�}�(�����h�� ���6&%	ǚ�w9�I� �WLNq�����)�Ħp:Q!?��v�d�FLr���5!�VX��o�v��MPy<.��#$F�	\E"��Z����g{#�� qz"�Uݨ�������5����X������=D��A25��{+J�.��P9�?�,���; ʼ��"zt�q�A	���5IK����)�i�!����]	:f�N׹�������PY��ln�5A�n.m�;:'ˆ���[&|E3\��Nayg����C�ʢ9
Z�K=�D�6����)#��(7<�ui~�h��	�XI�2<� O�Q�N����%I��1iz�@KG���!ۢ�딱Ͼ�~���ņ/sA,p�ڞ8�i�X�\��[���S�}p;}�LpB(Auk�Q���G�����\Wd
�%ɢ��|���56��bG�'�� �	�m�QAUS�2M�Pű#��`3����o�"5r��x�S�\1K�	�F2<�:���B�%���o%ho{o'"@rNM���������$3�Y����/�rЦ���=zi:'˝Ҿ���<Q�IkN֛��.����>��%/03����..���O[*Q����3��D)ȪfP�'�c�g\YA��77PH4���z�,�ņ��W��L.���M���G{�@�$�`��e@��~���r��xz>෠���v}��xC�{_E'���Y���@-U^���WD�5tf&-*�O���6\�50o֞�&pV�4߹4Ve*p㷦#މ�F�F.a�;�̿O�7C@F>ә�P�x�B���fV��i�����X)�IS���qLj�tM�ɑ0��#I�)��Ŭq)�����U�t  �=�ӊ��g�,|�}��c@nj��?�����%F����8�j_�~ �E��a���,\�M˷ Kkp�َ��N����v
:�N2���� '�!Sy�'[^f��d�"�O:�4��4���@�ïX�xQj����{"Wj�EH�i8�.��9,Mi
���_�J]�:����b�J��"²��w׵��
l@���t
��C=�d):��#6J4βI;�X@Ԡ%�wd-�*c�I���*��M���`$��WZ�h�+�}p}&�����a?�f�Xv�gW��b:����;!<�՜ȍY�ޮ
��0X����#=$��������?�4��R6N�B��@��h�>78�}T�I�y�α	-փ��F�Kj)�`a7;�PWE|�b����1��<�GQ����װv�+5��y��2/F��
�O;�?@q��u]?�,TP���l= ͝�/�,Ix�t�kCٞN�掉�8hB�s�m:"�fX��w{º]�dG�(
�;Q��0u<rZ	'��}��z�h�_H�D���\���K*�tW*�-�G!�%�ը�<���:LB���>?xkx�rO���X���=���N�1�2w_f����/�B�-�ż<�՜D�HGlEj;y�~�sw]hX<��T�?�џX̄�h�ƾ���g��n�	��}���QJl��}oݷ5�����=N՗@E�Vm�%!^�P0mc��f�)IҼ���H���BCk^�z���cKs=��:�����6��tjׯ������E<�y��:�Y?蒽�"ȱE1^o�����|-��a�=��M#�Kb�@%q�T�vR3��;��<fh+d"���#~u���o��|Di�B��c��E��-����z�(��Q8��j
�����d=���W �*��&�9$��/b�໫D	���1F��.����`_�����۫��/f��'^��wT<��b>�֤��ȃQ��df �'^[�iY��Uc�5�ġ�B��ma%�߉}�A�8�(Ո�xF��JIL�qbل������s����z01�����?�l�kRm o/�;1�,@��M6�	9���b7�Az����ʖ?5���6��h���?��+s!�I�o�Z-��R����Av��F!�s8�xT�֜S�U&��^����(ҠK�K ���
��_x�@��7��L�?���1S(V˿�n��3��]�ؖy�fj�X��i�d�r��,�^���V'b5LGc��	�r\e�xKN��^��0�1�v��ڲ�&���EQ���rZIx��懸CM&_�LC Pw���BF Jr�{����ܡ_�zefQ��4;�얘�_���t~ڀ��bG���vLG;u�r�(� �
t��L�:�.D��^�n�O�����Ձ�a��7�C�g�4h�e�����ס�Y�2)��Vb�ݪ�CNc�þ��9��{����_�xn1��+�1Ep���v��ּ�
��dr��H��ƭ;�*�MDN�1j �\�^���ݦB�x��,!lX��i$p�g�s�@�-	�_}f�����_a�Y�J!�%�Jf ����بm`Z���lq=`�8i�k2�4P���kߛa�<��ڱjڀ��M5ʳ,������u��	S�E;�ر�+o���Ut���Ģ�/�I8m���i�*A��,o/��dhŀ(�W�{�����R���H�L_�r�)"���N�Y�g�7��$1/���o�&� ��U���'U��7�M������YY+�Ǖ"YI�t#SqVNZ�Fv�FwZ��߆�p�!����?�o��*�o�ʝIj��DS��r��̉��-�H,N���M�FIK�=մ�w%���������D!wç&e�A�w��/l��$�T�{��A`E���$(񶑱"��[�!����@<�Lݓ,�(ixN���̂=���� ��'t��l܋�p���"���ƍ�K4��>U�׼6݋��B"��Fw��p9���r^����&�ш�SX/�-�D<ս.Y�G@�+˙��=_�$h�L�Ǯ��Җ������$�|�>�v�/@�!�9���������s�̝W<:����d�Ye'�rDK�A��.KF$<׹?��2�i#MCI2�^�}���;v��\b/��Ӫ]���g��&Z9��PA��� ;�ǂ�&=	,�Iq�F�����UN"D�
H^;Եl��5uTU"|����D������M�9�KI�t/�� m�D��,�؀�L�JX0��g�VB�RnU�JOt�L�S w������R��z�j��Ƣ�78m����ե{������~��a?�тa[����v�"Ӭ�%K���2}&֪�?�8,���n���8���<�Ru��W���	��C̅��B�Q��O�&��S�}��p�x��aa�`�q�� )�D�ڱ�}��X6�����t/�ͥ��
�	���R�5�=��`7��H��p\+�z���A���`���/�an_Ю�!��rx�lh�iu��~�bT깾QK˪x����{�����]b�kGr��_&m�'۲3�1��޽<�1l`�hu�qcm2}��E?�q�X�DIN7�Ǜ��;����`�{Xd5-c���M��t�rR`N.��S��R(��(b����P��~`s@5��">I@�������1��AU ^\�A���[�xȶv�Ml�T[Z�Jp���2�a��ӧ^Xv[-�?�r���'|��-,�1OP�}�M�d��ʾjf���RX�ǣ�X�L&�b�u~�K�.�	fytT�*��.tig����./���|�jZ�y�̮b�)�?�^�v�u�a5���[\%}>�״��6�P){� ]�:��}��_��Ƨ������m��"��
: �۝`����\��L�����mxAu��Uw��{/7ɳ�i�[��57���i��ވ��߇޶��5]�Y]�F-ԩ&���/P�:����/v��2O�~|U��'DH�2�]����ލ%��(�t)�i�ǰ?';;?qP{���:�w����fT���\x8���j'��ȍ�x��u�@g�Q��X8t����/�/�����l����-��)�8Gr�0�%5D�� Eb�>�2�(_-r`��Lە��[��Wp���FN5]0���e��QX�3a��B���P���j�o{t�^�;�j���᪤�J���{�q�����͏����s�P�۵ tH�6n�.)�n�HQ�`e2��)x?F'L>�\
����bI�g�RN��x�T����ѕ>#7�h�8%_�E�O��V=u7%�����y�19��ݵ�&	�V��Ä?�� �A��0�[���B�R�<���()�������ro@45�i>?C�K\=����~��׵�kƭ٪��;%i'��\��bx�5�W\h�ߏ����i�KM�u�u�}GtX���g�d��g(Sɮ��Ț˵2k�5�;��}ٲ�R.r�,
v�x!���5�C��-q,�6�yˑ ����/3Dx���� �}�x��Z�s�/�xn��O�o����Ns� �
np*(�<��%RԮ_tz7��H)`�����&�]�!V�dΛ�0~@��R<�(Y�q%^�A��s��8�f��fwZn�(���Z�N���v:\�9H�_���D�<i��~o�M��gM?����F�]��Z���%��P���WE�{	5�ݍ�o���v��T#��2����9���?�S�6�Ѵ�'��צX����K��0���3C�em�32����xs�5-����tq{BB�Uʕ�!E ��q�x^�����:٬%���G���C�������[bq�HaI���s'"��-��Ӳ��|!�A�ݜ��`
*K-L:]�u�s��ѥ������HO�KyC�MB,�I�F��_.����m�1kF �>�j�FDq(@^����;/�-�$!YB�i3UԻ�g��e���e�-/\xVV���v9!�߇��{�'T� ',l|o@��q���L �{���Ł+���B�����>shQ���'�$��||��na< ���КO�j7z-��Y�N闡U]]-p��V������G�G��vJ��lwr���k�M��6�<~��y�8Gl��j>K�שUz��5�9��p��Ds/��nH<T������ѣY�� �9ZT�	�gmU��Һn�+4�]�yV��1J�����p�VR^�4�����݂t��Ħ������U��uC7�u�@�#��kr$(9@�$[wu?P�LL��&('5^���C���&���R�A�Dċ��Ќ�Z���Z!�Dw�u�=�j��}�&كO�
ɫ�NT壘Y�%&���hTb�\�ް���6�+�I��䰧��$.x;����;���C.�p3�	.!�n�V4�������/�/1����� 7s���l�յ}��	b�rM���5H!qU�Ѿ+M`�1��{U��Ymv��4�ҍ���93s'��Aݚ�K]��	�ٺ%�� ���T(�`��{�/ȑ��#-�^��خ����tK��,� d8�[*�gp���*@��5�κ�<M{���z�I���2d����W0Ƹ_~�Dd[ �[�<57�.dtG7��T���ƃ-7h�K?cC4Ot���f�:�ow?�Zz�������d�������ί���̄���0��W~��f�����z��*߾�U��9�)�)x��w�F]C�Y&�UѢ�f�uP3�N���4���/Ɗ*��)��MA�a�0�E��W"���(+��)�lsq&L��B�3����Њ�n�g~pW��S��֘�c�U(��x��ě������ߢ��Z��r�2 ���*z�B̫��O�XW�~�T]o�SMP 	{��;v+�-��Q�4��f�.����0 =tk���>�������Vw��c�
\�Cq�٫�xu��3�3�
� 6|��QGȒ�n�c_bkM~��la�Ve�j�1�����m��@s  � ;��w$�[�TΟ�h��u�}#�T��J�	*�
	"�^u�c+�P��@�)E<�4C8ZK<Fh]�O��pUZ^J�j���ʖ������`6I3�,�(Z��j�&L	d�7E�_
��.'N ����"�_��`�K�PN�w�<���J s�`=΢:�w sM��||�C1:?��H�� �l7�s٩Iׅ<�D)�5l�g?�h��@=��}F��#���Kn�ND!FA�&��HX��=t'��zvdN��`�ᬼ*��K2!﵄`�ϻ��ز��i8��Lv�G+��9e����B�dC�܋(Y[ �����J�r��7��1���+K�Qf���8�0(g%��'֑E�.�i�94�(>[���u��Ȕx�1����PQ�؃��.`� �ޘ`�un�H�u$T�̟��Ҫb%*XFR`��TD�¥����2`�؝�xMxWƨ���7��"�(, 2H�?�7p�l�[�� �������n���� &ڌ�W����a��l�T�m���	XYڽ���)"U�e����:��X��d��E�>�h� �H}��jl)���o���u��\�տ)wl%�B�A�ܳ����
F�nx]������O��z_�%sz�k��Q�c�÷� so ����h?�(ކ�����&��7�l%햸�Ze6���M`U`P�m��'/Iz�|�����i=1�Ҁ����'
����t����W5�K�=Te����G �3$�i�����z����,�Kk\���ER?镔��\)GMƝd�W��m)ۂ�>P1��Ex�B�
��T���	�h1�,>��OnB:VOz�<��_�`�ڋ6�Lo��s0���UO��㺒������ݻ%�3_�N�z��c��p���M�(��i.���W�9=���]���7�ɫ�7!j�b��!&$8�;�@�炓�H�1�V8!�l�-0�����~[IsĈ�)>LU���FZ��[��y>.��D/y\( [0[X�ĺԅ	]d�?g���ks���6,dZ��Ol��3>���� km�.�_����gӑ���(��ޡ��]�׃�� ���)�K�B���@��=3uSH	;���I:>�^5hCt��
��@�Z�^B��9�u�U�?/-�B,
=	�	']���-A�k�ɍ��3��;C�W!';�����0�����\��I�&�W����f�e� 9�4?�@�(�5��4"�x���5����p�\��R���6�pҖ:ٚ}�{�5B�=�(�z��*(5�_�X(N%_n�2����X��Ng3�%^�f�易�]���.,�h��w3j֚v	�>=�NY�~����G�^��޿78���z_#�+�(B#�7�W ��}kRD������t�}5�Q��o2_�f?zN��h�O��Ad�����C�Ze�Ř��!���&�����@c�C�|"�i��lj�� ���|�>� ���M�$��F�x��Hs��灾�����bJì�Y5�ҫ�c0\�a�ǦQ�>�����f�2�hD毽����N�w��Z��v�Nb�1���B�1e:;�~7<�5_�[;*J1j
rQ��TM��l�3�jq��oK9�=;(��G�d�O-a�+@�C���u}��O����Z�`�C��:�n%��"���*rȵ:��Y?������R���ؒ)��8�U�jj�AȪP���ؘj�7,�6gI,��(|i������<n��f�^�}�B�!�M�'
>QF�����mp�����y���g��ި�(LT<:0��^��$���3��%����,d�N0�>L*��x�S�H$O�W'$=
DU�1c*,�QF�9������uX/@�N3Z�&��Q�S@R������b!2�c�mb2�a�m^s�.k��aq\�9m2:`�.��%JPpw$���G�Aɸ���(�m�*���+B��C.��m>HA��`�'F�l�TP�سX�Xg7ФP�@��Θ��B���R����fb��o�@�,�����|�c,��?�~������h�����W!��ӎ����?�cQw؃� ��Ӌ&�}���Ik� ��:��Q��|��WG�簀j��!B�L'l���lP�,�B�����j6+>��k����ü�%��!�<>K�7ȫ�ff���T�����f*���qI2�|읉y����S��8f�����N��zsf�h�
oS���0ok��p��Lu*qA���x�@,�w���M7T?��?�ME�8�
O�I�k�}�J�b7�؛�<&v1��4S�Y��j�6���x��݂��*
٪����ǀ�؅�k�v�dڻ��\Y�i��U�r�R'����"!�������}��,Ss^����=�r/���K�)
r�Z��ip��l�Z�)�GU�[�G�Ɵ@x�k`mND��<�Y��-~R"'��WV�k�:�a��7w���`�M�巽���ܫ��m�8�[��k�9�����En�&=^��7���*�*�a�Ms���齤"�p�wc�,��k;!M	`Es�[[in�'W����������BM��RL�~��>M+f��f�j�a�s�s��4�����pdn����Nj�md�q{�Ow"(�����/z����hC[I�UdBRm&ڭMX���o*E��|�׹c�7/���D��Olz5�n������␁�߱�{�S��(A��2J�/�e�;YbA���-���/E �F��(��|���kR �9>�Af�X>�������M���
?$Ġ2�к+*�R;��h��Q��ܜ���tS�zz?�w�[�x�@�=�]�?`�	<,�&�lׯ��7�g�`T���C`�`�����)\WԺ'�n����

��Y��klCk�z6�n�Iqh:3�&�K!�F�6��K჉��i���u�֌j���SV #}ʔ�v��L�̛�ޯ��Ŗ�؉�3@Q��͵ߩ��/NDQ>���\,8�@*k6�,�����@��<�u4	@JȑD\ԒR��	$cX�d�M�Bz��m����rP��񞲣$��Ey�@n����IL������G&ډ���K	�9;� R -�&jvv��폐:Մ�\~�5x�]H�5�i��J�[2�M+�3��������]�u��T��!����/5Z�R|���z\��,�K\Iq�a�Z�~�1�~qpCB)aA�HB��v�;�,^���-ջ�䐼xl�b����| ��}&�m����D�����\�>YfҚ8Bg3I:��R�+ؗ��D�BRrn����2�B���{g3A��C�9RЉq	ЖA�IX�x��0�"��W�+�k�w��+��/1Ԥ�h�<l�ѪW���D3Vaa�P_�V�-�$�A�!���[�#��6��U�: !�bYy �Fjw�|�K��Y%�_ͼ	�e�RSŏ���Et�=��TO�ȯ�z_��ݍ#�V�����S���كk��k�`�T\H{m�e�Y���n���J���y%�/۴���~��0%Z�96g%��?$:�*;�nxY�f�]� wr11X�e��hɆ���z
ł���[t��ۇ����B$oK�k������벲��А}�|� t-vQ��[&J´��
Ƈ�Y`-pX%���ח��L�d!Y�_+�U
��1�nJ�dp"���m�.�e>f ��	Mcu��s��DGvp�[�p�:B��N��/_��2��^H���`IPQ�=����ݺC�V)�����cE�r�YIK��f����8�ڃK��c!�ŷ��ϡ�	u��;K��P6�4���>q�X��ݼ�p��u|���--���=2$6o��*-�9HV�U+���G�{6��=�$|�W��J��hgL?��Y�٣��|�`�d� ��)ܳWЦn��C���*>ے<"2J}�=CS� ��3��2Ǘw�ah���P���*_ҡ5�� �ݯ"�d��?��mF4|8�e�5��R?Lq�5s�e�N__!�Z���Òu-��E�V�eL/A q���th
 �~�5AĆ�)���Ȍq�K
W(@?�k��-��%&bS�L���y��d0���f�ز�S�c
�����-���+L�B��h��JOR���� \���h9��T�o�w�q�|��2�5e���;'����M���Eu'K&s�*jO1�8�$��"��t�tݼ��/'�I��Jk-��TErt��}��n�/0�d�N�Ĩf��7��D��&p|9�\)��qK(�"���EmB�N�ǬyS_.rk��ת|N�������m,,�F'P�j��W�ҔҮ�q~\wz=�;���)U���xM��50),� .}�m�l	Τ���}��k7|V��"�Df�H��r�<n�+�*K�U�߃R�?7��i��|ų�#Si�,<�:���)�VQ☇(��cɋq ��u8���ݻ#F��1��UV<�����!b�FdDl�����,\�(��ũ1�=g G&<��ł���% /^��00 �	��\z�4'o7>ӗ��p� �S��
1�R?��M���U���װ�F恥17Ih�T���;���DFߡ7q�n0��[�f���d�qtJ�4����$�J`�덾���{�/P�s�(�1������8!��(�6�qa?S'��t�χρ
��5V�Ł��P�x�$�]�׉iIu�s7L�X�z'/㙺M�f��W?���=��1I���S ���DG	�AN{�{�m�0s�}�m8��R��gK������ճ�T���//U�pn�F+ 5��M�zF�-6D!k����;�Z�!oJ8򠯊J0/��,���p��0GPg�)W����c���p�<��WG��W�ɍ����j�@e=��B�-�ޢ�������q��=�+�a�Z��%�~W��.Ko'F��,�S3vok��fD���D��E�L���ㄜ����I�ᴚ�c�V��є7"�#��Mur���IV��h���v�`�s�$7L�2'4uN�4�]��j-�.����/��pN���=���B)Q�&P��m[(Ԯ̢�A�$O�Ჰ����T-H��"���%�Y��2}���F�3m��Z��L�J�bP�N�X/�%d��M.���n7->�VLh�{�j��cPH]�e�K96MD�x���`n\`�]G�N.7gǮීkÂ���d��؛2�$�]����eH��]����T�(X�<�B"<'�%���>���5q��iMq���7��H�Й�_I����;�����Q.��m�O瞀�ܧ�:F�$2ҕ?��.Ͱ¢�1�e(���7c�`��9�@}CY��S��Q��ݡ6m��͇��������6�/f�����fc�G�&O��pKM����8�l� K���7��'��|C�
H��}I�`��!fBf�9��M����(a�B���?��� a�O�>I�2O�P�G4"���f�c� )A��;��0p*�&��_Dc���oƴ�y]��x��'�㚄�P�x6 ���W4xW�q��v9��I�u&Ľ`H�+@��3��t=j�P�0����J?sh[�������fx�Co��\��O��o�1--�x,܋�M� ��T\���V5�q�z-u&;�o&�T�?,��/�N$����1Im�J3���(�Hp6P���'=��ע�Q�d�X�nnx�^g$��_�;�HO���������~l��"���C�G�r?�^\+yў�A�}(��ૂ�)�f�6��δid��^����hd4l����4�Q�aIw$��7ޣ/
�~���sMj�[}���%H��;��`�/�XE�%�S�2��q�"�	/�kT���P��3�$n��J��V��&�������N��0^|�;��S0&��q�3����1�+sSQ�OXq97��~��E�v+�rc�'��j�e�1^�1f�p��
���]�9��L|�Z.y�/������
e��\��%-:߂l�U1ޯ5�>��4��ѐ4��e?#_���>�Y��s~�w��S�g���>wY��fm�vR���ktLC)f�O��9:}���R�1�J��ǜwp�ߍz��=v�4�Ye�#�"(vU�^J_��$����^O�]�V�j��Del�~�'a�!|��*�/!У����!�������T�6�˰-
E�#^ɏ�-*����1��$���k�A��B��R��"�G`�T�;N�#��K��-G=�e��SJ
���c���@��w
�3r��m�M�v
Q|�r��M��3�f��]����
*�5�J��5�0�vg���5q�Qa�/
�����k��m�Ń�����5q3Z�O�f�b�Yl��)�؆�g�@rO�x���sr�^C��%�l�_멌�"#z�E�㇟Nd��:��m��0�������.��n���Km�44L*>�0
�n��cj"&������Cyn�~���ޱDc(|D��fY�9�
�FZ#}?3�t^Kq�򕢚%0��[%S|�u����r�D��N|���n�ٌ��6�&�:��r��x��G��
Jդ��0�!׊�Z�Ofz_7Ц��QY���֠@�)�6'l]͢��q��>!o��ܪ�설��5��z���hWiP�K1��s�"��b}��6��YŮ���e_c��)�U�16�(�)��d��]9��rl�k�P|V�� 8���A�8�k��#�N�3����"�E�{�&]e��J�UF_+�䗪~��~�k;��,Ķa���: �1?���D�����uK��_�T)T�����6p��Q�6-��e2� �;xH���e��>���U���_N�ɞ�tܛ���ֹ+Pd�9��cD� �����/~��@�E�J�AZtE�?Ix(o#/���w����|��]wD��{7<WPiW(L�-��E�F�~�� 0H=���ﾌ ڸ�W��uj�$wb�16'�L��<�M5m�`�\�ЁE|��au�DBI$�{�ȆS뺂[FN[�)��{.���i�a`�!�X�-��<��?����jW�����|M��-���IsoAWĥ�Xʲ
�w���c��x_TGތp�����,��5�� �\S22}*�|�ָs��$e�
�.D��).�E��x!�RIR�J����;�$#��iD��#�C�V~���Sd�ș�7�:���������?E\ä!���z��ǩo�8�8����k���"�/u4���	+ۥ�n�]� ^��J��W@ ��`T�xغK�㮖S;��#�nR%h VB�o��y��(*�߃���N���X�'dq0(��Ik�,,7S�EƊ ��pVƝd�Rֶ陸�U��ؗ���>��b����A���*�^���zYJ(�N�}�Zz�
��[>�V�����ش���D��^K�ގ���\�� v�=QI����f��y�<G&�����l�Ȱ�8��:T��j"�ϚP?�I[�/���.�&��a��ܹ���Q���P��?[����ঐ�'�����!���H@2��TP��]�U�t�wlԜ�_vzeF�C��6'JnX�S`���dR�jDOa���	����Ց+V^JmA��=>���O-a�� o"~$S����"ZE��x��0`�ѫ Jr��}1�@��C5�s�����W�*�Xil[�%��(f�`?��+9�7)9Q*���^���3r��e6��Z��A]�����n.1A��2�k�+�ۜA��~$��A��Z�bE 4�����Gk�C�SfF��&���J���+M�F��2C�S<��#fY44#yd�7��X���ruM�W�����;5� �\�4\6JV�Nnz�S;�g;�eb��P�xb���ʆ5�C�/>����WNc��t�"�b�
����������P�T������8}yhN�S�5�b�ΨGdi'S�3W@D%r T[�����4{9��X*��X��I�	y����Sp�J�������/���*��h�ʧ���j���k�ʯR2��Ȣ�6��Q!�E�����Mߩ�b8e:��R3��KՈ,z]�#���2%�5����k�3���Ե���T|���H;7�	��>��7�����^�Arfcl]��o ��7:h�:��]Ci��pn���7�ٲb��T4�� �e�s������n-�d��u]����:��U�a��[�Pۏ#�s�&c\�� �J!�-=1�v��o�2،�d5	ڪ�;������h���]�5��/O�zr�&<Ŧ���,��	%b�,�d�Ƈ4;k.�ږ�(s�T3&Ih1�n�/|�M}hW��:�{�Ks��y�T�]f�T�ɉ��|�~����i��Nz��<�cGO6�B:��сri��s&[d����B��9n�1��_T�u*Aw�%����$�ؙ��#���
\�N`��e����C�:b�ӎ̑H�y�7�LQCr�_z�R��g)4bH?�ٔ��ȽB�$�X00@N���8͢��%B"����H('ȶfd��n�4v�$-t�[Ƴ��3í��'��� J\��q��6�g�� /D����'��a��R��Pܻ��B�63�YG�1�؈m�,�5R;�����|1�j�S���������Ы����@�=8.���	�xn�MF��3� D���	wƸ��4�-~�"}�$�L�U�$��yD2�����;A��=����W���{=.��#|-���Z�:�^g� ��C���+���ׅ���-�)Ti���|[�C/���*#��Nk':��RWx!�=�Q�U>�d�6%���>��g?�+����x��mUKї�|��"T��cm�$��g��\�u���iB��Ĥ��}9Hk.����ӑ"������=����E���·�� ^3��S�8c�y��%�~6�=�/���k!��u��������o���Xp0�� ��I��7�U���	����:i�іN�.1vw�D�(�S*E���eeg\QǦ���0&�3o:.I%��l�Q�g��Xd�~�W� ��J4b��U�8�� ��i��x��*޾�>�-���$�lxe��'�)��%�3�u�)MG�<s�}�Ib�FO����@مk�6.n�x��a��D
�'��'	��c�K���:�]Á� �R�+���5�Ҹ���q=~҄����z�&V(G�d�Bz���4��謴
]���?b���<3_�� v����*�W��r9�xsXP��L�R�K����Kܻ�\u-�۔���"g�6,���Lbu���g
��Z_ٮ
��~�q���"���&g4���Z��"��a���pXk=9���J��y��&����-���&�S��c��\��p�J!���%GOg�R���dQ㷽P�f�K��Ĵ�f:��(ï& la�+���N�@�L��n?#G¶9y:>	��e筨�ہv�81h~Z�E`pb���1"`U4�v��yv��a&��k��jL�Y��Ȕ6k� /��1��>��H��cn�/*Du����Nt�ڧ����1�)Bj�6�C��ykӦ�S�Oc�8?�Y}%��}��ʖ�v _a���0<H��gk��v�Wk:s��ڭL��>WT��i+󱪡5n+�wp�[�I�w�xC!�֩��ILNN˔;4)2���i�����I�-�*�\�w$=�O��A���ע��)���#��M<��s}�W�Ԇ�/�X������p�}#|�c��U#���v�+�r�ˬ+�d���$�ըQ�C�f�.4�`_�-��o�ݞȠܹ?� �� t�䂆a-�C]�>��8��vf���X�������&`i��?�BѾ;#^|�z�S۞xg�)]�}���hKg��˰Ӫ�[n���N�.X��1ݍ�6�>l4<F
��H�w�Y�\�WEYdEh9�e�\��JC,x���W��:�:#٧Y��y肉�1S;&����>xg���v���b傍�cWy�7N#�]QdP�Jt7�_J^��qJ#��DA��O�CD�H�,����O{48.Y7�[��5v��;�j9�{2���ˮj,�PAϝ~�R�uZ�I��C��i���-�mO�+Kc|͆o�7�y�DhPG����:�p���`,|b9'�E)b1=���4v8��l��[X�H���h�ΕК��K�	�γ4a�cy'��fM{�)�9{�#U��}Q�?�_X\ia�e���,3l$6U��W�v
W0�r_A]��X�>�+�#��p�&��,#x�5����p��@�rv��/B	o�
��n��*�=��W���v��I�q�T��7\��(����l�	�H��#�"EW�rs����~�R����a$Rm��PT�x -����O�(���IU��$�Q'g�Y���6���t�f��J�v���c�{���˪.���X�g8��o�A`]+6d��XG��I����s����4ִv�v��f��J��gd �9�ف�Ņ<�Lv��
w�1j�T���٤v��sQ\���2�����@�精��F���OP���>sY��5I�/^D�Ү�L�[��4�Uy-x���xw�1�}�G��`�u���{t��D��Ce#b$ʗ�~�����P����&jAU�[0�IR�dEx��ɪ!�������V]&����E�İ��4i�[�N�"ANK���O�dE���^$�^��b�fp�K���o��KPj�� ��oF�<!&�ыU]ٚ������rIG������a����,:+a14���I����k����E��U9r)��j&<�< �F^�I<w<e�-�%��0������H?�u���{k����6����"4��uF:�?����.	|�*�8!�4��yY1���/ʓ(&�h������2�7��W�,y����EL9��t�z�jɻJM*n�>��5'['>j0>W�i~���:�����{_"��S������%��>�Y�w�$�LI
DgϩŦ��"C���0�Ph�aC[��}pH�.~ڳEq/��)XJ��w�6Y0��9EК:�����`Z����+�ګ��an�"��m���ϝ�3{��x��r2H�^��&U$�-�7����W��N!P��N���XSa��h!焟.t��;F��?�Y~��я�Ru�M�Fo/(�%��=��o�c��v8̼��m�V�RT����WZ�h��_�*��p,Yn��&�R�����l]�"b��E�4�e��=�|��
<u;�n'�EGu�M��VH6}�'[���(��k^�<9=� wN�V4�;ªj� ��_�zO)sc�,��3�`xgL`u��]{.�d�)iw+������+�L��df��٣�ǫ��};� +��J�wa���]8|)�����`LvP�����S�@���נQ�;U��6��5�'oc�����zu�H���U�+���u�oo��7�h��Y��@�i
�{�R ��}�Z��:�SS6��
1V�8��2_���(��KV����]���7�+�+I��S����B�>���C���F�=��mP|�la�E@���䠞�cU���y����"�5�Ɉ���6"�6N��T�m������(;��1Xw1�#��/�h�F�O��3�� �>�.	�r�W���9._�9܂��7��:��M��&�����n�i۝�W�hF���,�̵B$����a240�k!�`��iG��L<�@���b^2׾K�U��y�n4�3��į��/O�n/Ѩ! � ��,7�e>�N���\�����1I����ۑ��P�����-�]�j��N�x]p��^�������3KNHQ��6$���L2��`¾�ĺ���D��o<4+�/3�}%���@��{	��|����6eGP�o'�*&�zW�B��k��� ������q����Kl�,���ֻ1�7=A��%d7�~iɮ����>x�����w��[ 0l��vU{�W����;�(��Wq�'��=�Z<�pI��I�I��G&X �:��`��TV;��g^�������&D��Ëu�|�U`�/<�:}�����QRWU[&�-�P]l�Y��/�(��Qs���n[�W9��2�0�PH���W�f,N'N���$�M#��P 0���ʅq&V	J�~-o��"X�-���I����9���I�9u��VǕA�_X�ܦ=Hg��>�4�m⻆P�-v^��d��tonwl�{�^˱�8Rĳ�.��U�Og��wMơ��ژ��ғ�2h�͕�|���UH}5X)�9�D��C������LZ��p�-�������B�_��r�����c���hQ��D'E,	p9�Ooc�.Dk�0���t�+��(�Z��On�o9�߇���>uZ����<+��ւ4��>'ѧ�.)F�m3\l'�3�\!$�E�_W��g�)�0ޙ�.�܀qlPy�ڋ\Oz�"�uq��>��;)������2�^s� t�ڕ3�7���/|��X>���$4�t���Bٛ� ����P��$�Zۼa�g��e@���u�H��K���w<P��؟S�������>�|:򚒻ʕ �n�ɛ����*���4S�7�^F*J��/ﶚ4
A���j� �i�DOu(;0p�$�\���Wo�g��m����0${��b�<�R�2e����b���(�?&.�Շ#f��C(1���uj��[O�L�3��,��B����+)�t�*ٜ
��{> ����(NA�獲��'/�v(	s�dW�Tv�������ڕ$�����X|_9OZ�#!U�>-�Ů֣�ݾ1}D6�69���q_���%<��dFҺ�"#���sD�آu�-�$���&�Q�����L���z.��Nh��l����*�m�{�i\Q�����Y%�_ð�d��r,_?wg���_��%����D�Y'�%K;��k�=�i��q�拯��(%�a梙�a\�P���pD٪�-���8Ⱦ�Aǥ]�ҁ;*�{\�p^��L�����#XG�_��o�, ��r���ڨ��[{��q/�^O@�w�zK>���mq=�����a��vw<6�)�:p���ɝ{9�k��
x�Oy�N�.�׸�Mp�_AIʮ�]h]ܸ�錍 �u�ꆚ��E��C�f����ą�|�[����3_�6�(S�V��AҧB�����vF�R�Zb%7�e�&�V�6�߯�a.������#X��%��Wv���x���<��jE����װp��z�J�gv'�u�h��!�JWXh$�r��.p��.���<�N�>���׵�DZ̺�g�J�@o�\�d�����0u5�DzM�~�2��U{6l����L�l���n��Ln�6��(®WT`���q�{>̻R�>r�չ(�����&;Lyq_�x�W�Zy�O2�~u8�:���g��i�ڌ{�`	g�("�!� �o���O��kF��"ź�oւm��&�d$ʠ�ؓ�?\E��Rt�Es��K<:��G"�i9d�!f�q�j.���r�xd�$j��P�n�m����z^H�r�q�oS:F��
^�bY�,�J鵥d�9�^��R�������s*vĕ�F�+��ã����u}kP&YE|�~=;i��W<�$U����T���q�h�OA�7j�N)������)���¹f���I_t�Ӧ���o�ax�O���[si����&QEK0p��gӵ��R���B��)HJ�_�����i�H�R���vB��C���%��F���Hϥ�ٍ�r۝-�i��B<Aq_dey��d�F��3m0̉�g���1C�&��j�ڢQ��7/���x5V�W���dϳ	.�5���r�"��lҁ4���u�����[�&\�RZu�D�+1u��؄��(�d�oL\�@�m��|eI\�m�~��l��=+��e�����B����G A�FZ����?�!Z�^�	����B�;/ꑽb�k�E����ߒ d����,�u��d���`T�$�U�~����R��Z���pO��;����Mnu���#EW�D$.��@|�7�h	̄mw�ta^[�`,��6�`�Ey�|�~�s<�r6Ȫ�U-�Vh�=zo��rk��=%�6�׆*�1ge.�[�"�L��'��Jk��� �J1±z�*�<^��H�	(��K������Ϥ,<�Q��&�,���¡P-��V�9��ŝd庠�*�˃�j,ml/���
o��c��,m ��9蘎����s}�T״���@eݩ�c��Bc4��@P�fnWu���wj�T7�*lqlW���q��k	�C��e�a�%�@�vʮ�!�B���7�~\J]	't��E�b+�}��|.v@��������w��&PQӘ�J���"���c3*ܾؽ��|��9�1 gui���ﵷ	��.qJ&`-��?�mHt�6d�Dr�6�d��F!YF�sb��B�e��@��=h?��"������~��~7lŋ$�$;������ٔJs0*��N �[�Lu���H0��a�ܾ�nʿ��S�m�T��F��#׷�!��Lɯ�*yҒ�Ɵ!������[�8�1	��X� ���?��\�Sq7WYUUu=�ޙ��� ��-�i�q��ʭ���(��|��g|� ��4���)=���G#u�	�Sv]��ʇbDg��]~��ҹ9�%vw�@��]�;�T��q3�H���� 4Ҧ��e�8������V���%�qD��&r��;�[��ɤ@��P%�L����r��v�����_d>/��h- bw�!R;�4L�FG
���G�(B�/I@���E"�&oӴ	�:��|	�k�F*Մ��U�+�Xy-bΕښ�fIq���t��XT�I�U�[�]�D�C�"��95-��䄔�93>�@Ǚ@��rɱ�I�����5�I��ja�IRK�8jC��E�Xx����5IK4XvTl��6F���D)e�1�{��@}U�T�������C�_e�y[�L�Im<�:`ag�c*'�i����k�^~��D��N�MrϺ�÷;�����홷��y�q��Gj�Z�� � |�Ã�yЇb��%.#�[�k	���q
�aҧ����e��]�!�yS�+9n�jB5�4��ZvB$���(|�u�Y!����s�p����֙8�uF-[�S@����������E��:R��I��!Ź~~��=%�)ݚ��q�KO9����l]d��3]��i��ŧU��'&��8�9L�!k��qA
U\z��G�v'����t�I��cUM ��D�Ejy��R�g�9ʘ�a>2��8W�_T�ogÚP邷����k���W�{6��oS�J׍\�[�g��tBCB���2��@,�@d�;�fo�;��}�u���jRΗ��"_��W�P��ƛPCѬB����Q�Ejb����+��DR ��`����3�~��*�=�9��0#��i�i�2M牴��X�Y6���[-h�1f^R��Zy�|tƋ�l���P*o�u�+���k��\*��*uv���Ȁ�4�1�Z�2���c���E:8�*p�."˕ݒU�hfÿS��Xz����i������@�X��Ѓ����}'�4��'�Q@S�~1]�V)U�� �
֖�K\�
df�Q�:(�2�����啘9�m�C��iB�\�{�<��T�A�m�)��:%uNw��('���`zO�����+�&��+�)��+J�/_����͙���H��g��	Z��/ju[��x*��\e�Q��m�a���Mj���-ߚ�����D4�ʞ>�Ƴ��CZ��0�~Z��ޫy�t/��n���C�� 7���0#\���N=���ED��Jv���:�U�O0d�N����r��x�JF�)�����2��$���ޒ�DZa�㮫��
G���a�����
XVR�v�G�P�y�u�<&�����C(r�tGd����	�q�8��I�p1�YԢ�U���d^��?�a�Y�k�\���C3����%�� Qm�����/A*�<R��`�t֘��Y�3or���q']LV�pï����U�26��W|�B==V����t�[��NqN�$*WZ�f��[����`ɫ��x����C3ezY�y���0g���E%��B3%e���.}�{6��G,y$����[�H��L>���1a�@�3
�ީ�ƒ����н��Ω�ئdwS�����AY��8����~�8����.��5�k���,_ꦎY��?'ջ�\��2)�\�\B&+k�� ��!ȎG�13۾�nslr�@����G:4�C�M5XH�%S���Q�{i��]\�H ��������}�nFk.S�	0�H\%_4j��k���#��B��𡸘}}��Wk V��o!貗�߯��ķBr�� Z:�=�A������W�	��.��ˮ��c�O��gX��]�B}�p�3BV����[�Z<�<���!�1I��:��N�cMk�'�`h�ř���?�{�R[�<�[�PԄTY�5T�����Cɺ������@WY*�y�Z��2�⼜߉C�a�����A��Z?ZH�b��%�םY�� B��ƞ�"0�9�@0{�t�ӛ��v[4��`��f����GĔ�8�?�PSN�����y��Y�n��T�jhB�[ےm��qRI�=��=��Ƴ;�UӃ��7#17h�-g֖z����� ���^y��{���?�<ϕ}c{Q������#�~�?�y6�7�Vtc}T�nH�׃��%k���,�U#A|t֋�z_��}3�rJ�3�H� �9��Ir��,��,;�&(w�B�ѓ�kO�$�s�3��G�a�{�ӁcE)U�����VC��]b������J�9:+U�Z�+��si��ZwqoY���j����$���V�W{��P��K`72��� ��r������ݵ~�/'�8O��3)�1���s;*O��ʵ����)�C�	�>^н��]еo�5G^�a�j�9Ti��r8 ������'O�Ƭ d������6gxD�f'�S���Q�s��7E�<)�yd�v<���iV*ll��WHfB��Y���Sc�	�ug/0-n�Ϫ���u�4J,} $�>�v$j�>�qXWp/pW���G{�D@����^I���x���h�����k����(&�����a�z ��J����^i�@�<{�=�VF��.��@�Yg_�����p�O�"�M�6��:}* (���W9a �渏G�-J_��(�a0#�l�Y�o&�TA��D�S���������v���J��5]�ϯ�B�H9�]tlQ�-�ZF����ݓ����+
�G���%�2�T	5@4���K(,v���>��-ٓ1g�73�	F�K�E%BO���=�|����$���*O+ncy�[
�h�#r�����ʆ�m/X����4�R=m�m�e����*��H{��Q!]�P�@���%���J3jDɺ�=✠���!��S �g6l�-K���B�E�;�L�z��������.��� �:,A�C~�Vt�9��,��JI�m{�JU�}��<n��}�)
�	��$u,/�¡K���xq�Y38m�w<Q�!��c�y�Qm�����H�k�,!hĽY�~P뺓�Dk�x-yV䬱#�
�隍�"Cnn��:�/���.�Md#@�&*��o\E'��6�hq��g�YZ�ױ���çX+���B��19E=���o�|iy�xa�wjo�)�G~�iV�ǏS���ƈ�1�^WZ�y�P�6��aVJ��H�7�:Y�<�nWs�X?����MP�@w禦����Y�W�5%��"���>��V7���K�p̀!�Ն�`|�"E������Ot���.Gy�!��$�3�ǋ�����봧)k���(����1�� Ho�Cd�B>.���N���5&�㎡���[$Bo|o��P���Hm��N�WWOg�FT��d�	�3��%g;]q>S��$��◹����ab��؈�͒N����xz�o2�l�d��D;�y�4�6J-Z���Z�u�n4�]V��ͳz�Qc�L6�a�]
 �`R�:��G���e؋�hl��@�?�-��P�ES�Z�S�j������$Y7%<CV�V� ����sj����'�NU����c�4���D���p48�D(�W��@F�㤄8]��#�TI����)�$�#��$��u|����M������Js��Q��U�ҳ/ŷ�N�ũz�����^w�k�D���Q�b��#�t�= Ja��'������VL�r�����͚:T����(!�^�;�� �W0��m�P�:_��#��:Pp��sZ,�K�-K��vљ3x��}�UEBPn�_��R<��a\��]�p�z�
?$Ry��F��D�{F��E�1��E~ҋa���+%~r�����YG��*��Un�WX�\������*��_�%�Y~l��m��pJN���E;������H�ܫ
x�����づ�nqV��,B��XA��ޝ�� �>�� vQ��qX��Z��s� [x��nk��)1�ڀR)H��R(ՔX1�/K�E|���]�$v�,b�_I�){Ƨc�C�i�[�9薃!ǹ\�U�(*�`@��@Qܲ����=�'��p�!��h��''5��aނ�§�2�v�F����E���Yڨ�P7�-�Qt�v��2};�Ĩky�������zy)�[oq�.��2�c��:���[�LDn\ᅨj,7d���RE_��� 8q)�]3��=e�m�*�\@�{�]�P;���asц�c��As���g�	Y���3 �_zY#��
HJ��eտ�gyv�H(֋�h���z�X?�d?%�բsI.^hH�J2�ȕ��}�a �V>�7�B�c<��[s���i���2���NoԎӨs4(/��x�K�(�'�?�0~'Oz������
|�	��C������B��Y��58���C�R���L������[����������,l-�I٭qd���Q3��Pa�|af(���5��;��E �yJeR}�;��&�쨣Y���5�|_�9N�X��2��:-<ዊDxt�}���,@�uX%v�C�_L�$ҥ�7<g\D4X��4j)�$�Dڊf1ǝWp''��4���Zr��Y^z��d=%���hWWӞ5��5�{��o���;��Ʉ������#����H&�г�%"��f=��1��Y�R/cE�n�UϽ����/Y�	XIt@%�H�����aQ��{%(��QcPcڗ�h�}�^�@W���1�AYL�?P���E�l���ؕC�K��+xC��< �)�f���*pX�o�������̉y85(ܐ��5�g�ֶ�Y�
��cJx�Aܢ]��y�sz��}yf�@{�}�I��3�ߒ�+�WoH�'Ӆ�m�J�J�'Ji\}>7�0Mܵ�Ia
n7�H���Uꓸ4	�����5�o6��ra�O ��hz��Vbj2�뢵H�@�]� ��$yh�������5��6���� ��>���('gs�)"��ޔ1e�Q��:N�J�<�YO\1��X�%��wV��c���-��Լs����k�R��|%](��Up�������j���T���/��rB��j�4&�'p�/Pw{G �j�t�Xi�љ�d<~Hp��ǫ^�L�C|�{�GP�e��:>o,u��~���mҧ1�)f0M����/A��@K�Y��?9�b��i
�3�n�dP�'������]?~˚iL�Q��(1D�tD���)�|g{��UG��r�^�q��@}xLO��TuK�#�}ChT=C@>��z1(^�j�1hS��gw9�������j@��n�4�V�k��T:����-7��x:�4���V�]k��2�h�S*( nX�H�Ӷ���A�~�fa;��, 	'tq�����C���?�m=a�������AC�A���� LZ�4B�O�Z�3{��Vį)E��H�u��s<a2������	#��K�%���8�YH�/��'(�?�"����� �l� ���T���"v�p���'�.hΌ$��৐��`A9��׼���v��s���|>]f������=��4l Tt�I�CWd����9��l��v �o=�E��uX�m�)$��5+����t��.��D1��W-g���R��`�%�Q*��^�B�C[3f"�e��@��յ#��0�A��](�M΀��Q��	�6= x�w8U�n���Hǂ-V�)��b�>*��ЅM����U>��) �*�ܧlЄ�<�!sJ��Vj�o���2G�G��K��a�A��ç�W���+���ާu�%\0A�yZ�.j-��� ���.���E�֭(�梅�=�.�}�Gf�:)yyN.3��\�w�~q��m^D��;��W��5�?
,Lt�ju���T�Χ�;CF7�=*%h�u�7��{���ָغ^6�A!��ā�ӄDo<����.��qyu	w%�Km��ʿ�
���j��皜o\D�;7��}��=���8B #]ޝ(���,�����ô�N� ��T=U�;����{WIls-�9���-��RP�� k[2a�z�T�5R���F@��] =��2�d�'4.��1_���*&����͂a�-������� ���X�nyQ>jl��}crM���@}�d�D[z̙�H/��2��c�I�cΰ���	�׊��g6N�=Xe>�3�/��@;?����9R�{~V1K-z��l��GSup�2X+X_~���I1}�_FFz����\հS[�-��^�ˍ�X*UŖ� ��Z�L�`Ve
C"��h��:��˔pl�Z!_�rT6�ښ�
��U�jh(l�r�2���_U��*���b�ƪq��휮���鳜H�����dՄD|�[ ���׭����,t9�F)�j�gjuU&p߉m7/�٢�v��|��4=KͶ�}���;��H��O�R45A���i�\�K!��'�$� �9��w(���榋k�I!m�o���nW�U�$�"(�Vq����[h�GM��,8�#-�+�PM�)��\���7����S�*I:POL2�,d{I��"(�q��<�ς�A�a=�;��>�����:�0uʍ�cdg��_o��UT4�Ț'� |K�rΘi�O[���z-�`&@��@��y�G�ы)��s?��@��PJoΏ+N�#1�HT$�2�T��-�
�]Q���һjXW�M��!p�Aa܌���%��a$֕|g�#�M���و�1�'���/�^�F��>�b�=��q%"�@L-�6���d���E���TN���@�?��ɹ�S��X�}9$�boPoLᬯ��N����V1�\�R;�u�	E���=���J��"&eG��bL�yr3/�ܶ,|L!��d�i�c)]	Ё��,�*hPy����M����km���1��d�{� @� QS�8�y��/ɭ��pY�KR���rh������(^uf�?A�ma&��(�T௎���pY��ʂ
�����aCx�C�u彜o�b,�k�̮�~�j�J6�P�מ0ӵɑ6�S���su!Jf!F����Ii������O*r�������ˈ&fا�^��7�2����
 ���K��"*\Ǘ>�9�eγM��5�1u�4�p/��/�,��{Ǔ��۷#"���	������ ���.2��[
0�$�m�v\!����w�gFs�T\��|��"�P�'����<��[�I�t�Ħ�&z���;o)�\���½�c�=�K�z��`�CJX����uB�onP�<K<�l���CnDv�dT�:j���R�}�+�T�E.�Z�Cnf��©aI�&�����F�F�.KS���k�j�AwƇ|^;,���t�zk2� ���� ����@D�a�����q����{�X+[���-�\[�qr��;������s���rɃt:D ��������+��	B(��h���>v	����b��W���z ����I���ϱ��n�$P��5�x��H�ȃ��d@�a����ѭ:�o���^�Ϳ����qVT���S9ߍ�S��n��v��!��'���j�(����M6e�k1�S{���H�_�]UU�]Ȳy�� 0>�0���{#��/�?$��E�W�Q~��P?B.��F����\�U�g@�Z��B�X�;g\���;c�U�f���5�x�,�jR���X|�B7����On�-,�h�W��K�QAS��d�i�5�Y����0>�Fx��e<rp0Z1̢�]z�CS�7}�%�)�	�e��q��u���������r��f.LԶ�A�� ͟^�l$ഓ.�`eo�� �̏C�W��b��
�5� ��M������`�&o�D�>o�/�L�1��|���rn������nA_L�,�&���䲸@����_A���׶��q\`�R���A�ܪ�`�R,2�.M���O����0�E�0���.�C�Iu%�=�����p�E��Z:�����w���W�4��n�=�����u}�sh��	����X3X�LsRv��
��	�8
���	�x�&�t��c��<`�����Wg�͸�1�M�>~G9`D8������K�S��M���hg�ا��R��#r��(���e�_�Z�&�
=E�-w���1���ʋ!!4B���zؽ�s$f��
��7�{s�-�P��.Qo(��z�p�&���&�@:ҋ����[�����zB���������Q���f��ޱ;��̈g�޿V��̏���� ��� 踘�$�&�U��!("ͮ$�q�8��	FR�����'C�c���0�M�U1�(1�ܴ'S�1��5����T�{��lIL�\�N:�k3�9L1�� Up�T��Ig4D��3�:�s;r��訨5�Ki"#��S.�>���}�����6�G��j,��ېq�£_��M4u�H�@.��?�B��'���T�u�������A��{YMq� �� ������C�36Jɂ��X�'�ľ?rv��Y�#��
�I�i-bt�_��lS��q��TI{���\臶6
�V�y�c X��P6Y ON����s��d6�@�O v��(4���j���i�]�z��8R�1*�ʚ[R�_Ǆ�Un%�R+�\��|�����t�h=dz�,#����1�������Gd�x-��~ �F�x���Mz�������iT�E�6)j����P�<��+J��߳m:�u���5�r�v�*b����p��7����e���q��K!��UT�-ut�Da8���v���Jxrv�窏L@�DA��]���I��;)F���h��r�('��tVܣ�����.oUb` =L
z�x�L�gDV�/.F���(o���= ����le����x"����� j����r��F��77�O��A��`�,*�pΪ�*!KJc�O�uء��d�)�`�轙���%��5��+��!/�Rt 1�� ˑ�T��Å���
,�`� 
��?�{ɔ(�般�7"��5V˱����Y�o ���T���b#E�G�Z>�Ų�ݺ����@@�@�5h.�Xc�mQ����힔$�e`;JD�įp#�8h�4M=#�5��v�]Зs'�`�d^}�:��}��BT�"�$ڞ���(AjUl���r9�y��`�t�Q�ߢ	�9 �U���+f8B�ZւPl=lb���s�Sk�݆���
��%���{�f���i1����ą��џh���V �ӷx!���|��辎��llm��a�I-38�J�B��_x5��aB��F�]c �ڷ
���m��p\"�!z:�x[�U��Ǣ���Cֻ�r�2�F�E��(<x��;�ɧ'-��SNJ�o'���[�|hi$⡍?�t����s}�Ҏ�S:��Y�6�j\�y�ӌ�vz,BVR���L`$Z�Lbn��I���\�5��j�AXz1���e �%�}!IĲ��F�HEȋ��	)�&�h�J�֑m��v䄬�p�깩(o4t<��G7��ZI�=a�}�,tKR�yL�>r!��H�Nu�f�J@�����뛘z��O��X`�9�8dM���ۉ~lr�r�v���Ë���5��[�]���h�[̸�1�3M�rG+�
A��;���V�V�5��i�Q�sx�����@��(⩭|5��[��Uw�of/���G�� l���M��v\���AP�.ӅfL�̆HǪnT!���k�a65MpȠD'�*%pp%>q/܅)!$�o$ل^�n�1���$ap:ŀq�[� ��� ��ғ��?>���=�Y)lP���@]:�oj���N�뾞�(��.$A�Q��S���[�T ;e�2/}����!m)�2^�}�.��X��Jzv�򪭮_z��дA�A�y��<Rqx[9q�ݸ���\�� �E�t�dx���s�3�  [g��` 31+�(����v� � ������I�������������W�l��jJ�8e.�eT) J����"y�h�"�+���N�[7�D�>�Y�#�Oh��+
a��'t��*6aiL���SA�I
O�*�A"�G��ed�;�+8�j>��\����Y���D�o*���s#�E7�!i���}�ި����F�C�"G��&�^SQ]�V.�uK��҇$<�������Ϗ� Q!_#r |�	��m���7����Ř�:B��5TӨ�G?��kآ_��:��+���0�*z�V��A�<����W�2�;�� �m�i?AU�E��4O�@Mq�4��nUu��y�Y��IS^ Y�i���eQdՔ�CSE��s�`��tLB3��rxS�B��<���Y��׳�u�]px�j\W�+�P/�(v���X�Fg��a���y�ތ����Ӗ���;�q�0��嵳�pH��̶��z�,+�����}���mg+q�.ז6�;��B��?`�9s�4��51�(�����j�"��g<��yܻ�쇯�_rs_��R	�2OFYgT,�[e�<�b���P���9m3z����+�ތU��F��xvX��Il�4����U�L`�dP���w��EQ���
�)R���v���T.��"c�"�H�??�M��~�3�KW��� P?ۢ�$�bW�N6;utjp?��a�mxE�o{�0<��D~Y䱦�w8b"���&?���I/��:�K
ƌ�u����aa�:�W�o�j7�+�Ϻ�~�� ިN��B'�]�W&��]}l���OZ�� w1ǼeO��|f��|�i�&����H��	��jy��d@�/�� GD!�
3�����Bk;%�7;ނ��[����h�|�U�q�u����+_�2��������$��pKF��Kս����[ynÂ��}�a���C��[�+Ė�e[���S��k�z4x�<֨��I���*|�ͱ&�9,�ff@�(�LM�~�8�=;3s3�K!��5qf]o��'_ܩn�pA�#��G��d�A����8��HIY��U)��ؾ�� $�����zA�������#��0L.̯LVɻ����Ҝ��C_ͪ��/�yL)T^⏥�)�5�[���Z�V�n��6ċb]�Xŀ���2�4���NA����?�#��U*���.럜�,MA��_`���'�P��ՐF��L��?�h��R,|��@���`)f�����Ƃ:<Bl-��ûu��z�we���,j��4Қ�vxۮ��ro8�؞����'똞΍��K<�J9Y��W�*����]%GrW={,~y'�bW#`u�B��4-�^��Ƭ�<��|����2IS�[5Fro��+���&E?�c��I���*	U�kY�ݝ/Z+�z̊�< ��q�6��TL\(,���_��`u���C�e?�;c�V~�Y��b&���IK��7	���O�� ʭ�J�`x�*��P�I�4`��k�O���V����Kqk\����Y����e߫Ǐ�=Nv�j����#����@�4��tu�_Gh�$�ox�?F5�V ��p��G)Z��L��ND����Q-֔�)���8^?`u�{��/g.�3W�P��)|M%2�"��]N�g�l2<_�d�9`74�y8�QlI�� ].B�
#
�i�g��`�}o���t�dA?D��R����fŶ���#�:$-w�����H��f_��˿��;��馈�9��{IB�όQ����E6�2wx����9�p�3'���4r=u�F4wU����$x-�P�D@���,O-"dV�+�]�� �-zM�q�A�����"���"�� ��O�5vؿU^�eJqc$�w㑼�{4�~����t�^ccUI�L��p�*\����g�~M�rT}��#�o�i�T�y ��������p����FS1��E�x��?��.uʚNj��$JՂ)�a�4b�3|�*�ٗܩӼ��>�#��Od>��O�8��xu�fŘtB9ͣ>�<�np��ޤM�70��r��?���WӦ�Ķ]/%P�l�r3�K9�J�_�հۿ�ߣ��k�tX�%+m@:Yn�K�c�=��b��kU�ykR�*G�K���Q�\5S�������7�9���3 3�ᶖ�{��̠観��Y�R����@��H��#��H9~����{�YO���X��Zy��n�g�Ql�?/'���3�`��k���(d�Y�����Q5�@���h� 3� 複�>{A�r�ѮGO��,�, �Bg��e��Ϫ�N���r�V��r7&�mQX��PDK6�r߈�^zT�Zd_��U[��=x���'P�_��c�K%q���	�����l)��\����i׎X�U .�'�u\c��\�����2������AF#҄�j��+SgU�0I���B!�FJ�fY���n�fY'�G��JN�+�|;�$)�8X���Mgw�#��%sW�A��{=�8��~��>�#+&�	l�<���{����N�5*]��}�*��l-ޔ-�L8ە� �N�13'T�]��f���U��}���27�OG�_|x-|�0��}#��˰d=!`$)����>�Kk&A�� ���!��Z0�Rdu�� ���$Y]�$�U���y���0!�1߶�ܘ�י;��3�[�EC�O�P�ۭpnݿ�?�;��@,4`S(��{�DKàm�Ҍs�l'����J�z;���]��-���
x`dQ7+�q��?��Y��Q0�o���Bf
?ٴ\�R'� �#}^Gt�F�j�c� �UQa�Ad<�������ݡ����|�\u�~�jx�N���h�y|�ҧ��f96���5���|k��N
ZDb��蘿�� e���E�5�ǂ�[�GA9Z��qR&39J��Z$Y�E+X�2�ܝ�Y(��»帠����R)�*��w�sw�>ց���d�љac��:�.0X�Q�b)�k1}����F�gm���d����Eӏj�85���_(~̿��ckW3m,��w�G�J/�s%ؤ�9S��T�t������}2������=Ѩ�py� EY5�����(�w-��~l��=�|�=�\(��I���V|DX,�];�'�U��Q��'�t��L�ϛz	 ��{��43�w���S�5LhY*��=[q��ަ<Y;}bCtH�_D���jPNv���CVt��f؊_�j�>">��fʢ`#K�c��g�γ�t�*3�����;W�w&��uQ����a��t8'V)�%Ķ�U?��]/+�@�'��о�@%�Ё8�^	����g�l_�|s��� ��Y�|�A�4�<��F�CAHg �O�V#:?q:s�_.#�T�;�.a-}�G���>���j��VɓA} ���8�'�=�v�%�L^"�&9W}Ϩ"
GN�7.���6�/��3^~@�!,z^��¶|�}�8�f��KF��q�7k�������*��J�-B!��v������+��k��n�)n�L(�?��̕f��L>F��C^!�>\X?���������տ�ND��)f�+'����0%&U]��c�����{�)�����S�� 9R�P� �䪕w�t5!��b i@�͓�	y_�}c�JBNM7���EA�N)j;��u�D�?7L�u���{�q��ld]�G,9X�|��3������u�a6-FS<��8_OF�!>�����o�D*�cZ;<΍mYg�Jsk&P��vUE��h�����$�(�»}R���[�/0Sp�N�=�=�C-��k�1{]�X' ��ڡ�ŋ�8�v5��DIWX}v 5B
i��N���=�|*GX�9��������l�?���ֱ��d�����Կ����9Zp�nϧ��0!�)����Վ�����c�a	&&Y��e^AQ��p�~�_��T�L��pg ��7�52�u�`�#�!��φ
���Z	�]���'a� ����=����u#^���ui5oNl~Ke6:�v��^��H��7��;|_� �Y^��_5���r�D�N�����y���:��/��;��{y�\m�M�b#��v���r�A��N�R �c�-�d5�u�ZHQ_U�,�=~B��>����ҟ&&��y�b�D���q���U ��kG*��=�P�tB�R��V��H�dG�ף�2���~�@��k�hv̘�j�1+�U��k� ��L�p����Xmc��<�B1�~ruC�o���O��"�H��9�V����h�'���rc��`������GXay1U
L�T�(R�5bvxA���E����7������ �����3�����-��b޷o��+���W�%*�0~� �*XZ8�d��d|���{�!�
�O��U��4��E2�/�2�eҾiA���P�3�j���5M��UR*���-�f�x�T�U�L��(Odݷ�zCJ�d�y�PL 
h�h������	f�����N�4YS��1{�TM�W҇�ι7�qO�͛U��x_+' �M�"戄�o��[�P�0YX�t����+]���kW�ɲr&l��Ԓ5;��l`��0}���՚����@}*�s
����<����i�] ���hI��}�3{��KS��=���:��4_��ǫ��/��T�P�S�D�׈L�;�%�B�1;/�/A�ԭ� ̼{UՍ�ax4���._ ?���4��gf5�$-��B�����Xz�ѧR�r�Brs�(y�~2R%^c7p�@]7&-�n��՘o�כ#�X
f�W׳Z���4���|C�B3:
��;9�(o�l�RKƵ`�	�@i�`��.85�FM4�:%iKi7�{y_�oH��H��@�Qr���|ؚ@ԣO462 C��m?'[������,��X,�~w���|�@0)cm)�ש���q1.ǞIg:=S��4(а?t�\�b��k��G�̈��L׈���f$j�_���j���w��2��/���f��w����8*N�Fa�OW�Eg���� �%���Кs��hO&�~�ۊ{�ԭ��z&�7]�;9�E��r�Q����y���G"짟�RI%�*�=���蝸(��N�=&��a�4�O���YO��ar�u�%Qj��&�*"��~��&��g+ˆ�W1z�[oJ�͛����"�-X59�{�d�JT��/ל�r���K�i#�����-t��Ag��9��!��o��yǨ���)�������p�c�F��WUtg��>J�C?�m�.��]�'�sތt�K2���ܲ,���>��"MW���=فH�,����a�����	?��p[9H0=�c�=�ϩ��9�n7/�L6�w@���,����a�rB b���
I�0��H�w]�AsS�8����ٳF#K5w����Y��J�K��Y);@?��xnO}E~xj�{U���6n��)e�^Ͱ/ty�J���X����n�/�3���>�rgҍ���ml;�7��4��G6Νt�'3��N���l매I�t��S�|��vF���>�T�rx�Ő��Kԁ�� *g�n���}x�y����Gj�8-[T�h6G������{J��G8`G`$��7���N��'��Y��PS�}��(����[���p��otJ��oۻ߹�[C�"d�*&.�y��V��~9���<�c�B�/Cx��4�2�&7_�^�S��i	�a�HQɐU�'��xL�XL��9V����g N��z�&u��^�C3oi���I �! �JgX���y ��p��8.�\����:=h�`��M�]�(��&Y�s(u \oIǷ�����H���:�����e<�O�L�M�]����o���{l���;��k�ւ���c��A�*�7�!�y؈���IX��;B]�'^2�Z,�� �޾+^�0zyr�����A��yo@��2J��I�''#�s�7�x��x�'�:Xء�4��\X��8�Q����-���U4��H��%�2wvr�'�)�e��5y��ތ���R���R�L��]�+P�md,�3z����yq��W�۷�rL髅~0�,����pl�sJ�FH�VRU���=t��ϐ������E3��A�X���:��������!�=�*yI�7���kR΂����=k�0�"�s�#��X�j�#��G�w)��>�So������l�lA���5�Y�}dǗ
r�Ň�bb���#B�h���=|[J��UZ"�p2�+\�H�	7jP��%��Ȏ�Y���`�/mp7�r{]��
7m[�"֚$!��"ΔN�L|i;4���2��:v'���`W9\�^T��r&��v\<���B��0��������ϟ�}ʻ�Z�����i�K���u|/����]s]i��R�ql�ލ7ȹ`�����v���IXB��v^�W ��CS ��K�(6�	�������/��hF�󧘝@���q ���-؉#r��������]n���Y�V4����E
�x�E;>j�T������� �r]�����ھ�Y��:�b�C�G�*I�%��2!�#��;�.91�T�f�bp('��&@?Z��A_֙ܖ�g���JT�	��m�.������>����2�{����%̸�%i���*�y�Y}Zo�L���j�Xz�+�in�N��|.ݤ8�s�w�}Lh��d��R����d+Tm�����Ϟ7�L��K�u^��1���
�Muu�h��`<y	��x�H^�b���tI�"�Ӷ�A9t�8 6���r��
y��1�5�j@�~;�ui)Gh�H?%��HGkI�~���6�/�W�b���3��?�,��Z���/�"*��S���%J�r��u�#�`�����b�f�v���4	�3�Z���n/\9G���n�"���P��,/���v���J �f�;y�	J���f:����&(=�HAZ�^�����VK�0�fX���r#Ř�5`nQ#�����L�^��O
�1�_w>o��VG�_�4`�"���k#��|�XA�+�$�0w٬q����A|T@G�s��LMG��F��Oj?��+o����a<�c&WYN���ؔ���Hvm_�����R�Q��%�+]杍�W�t ]��@�l�PB�O�s�a�pz2�[i�K!�7����Y2pI��[���qS��5��A���h/��v��Cr�R=�bQQT1��� ��ξ�aB�i>"��}���j���̖R�$B�JXǳ�)���UT�I0r�,p���$��������O}�%�#���?w����w(�IuxBb!Z�<ߚ����ڦ-cN��%z�l��	�@b�:� B�j}z��� ����QM�+\.|��ܵ�\�p���6�Lu��5�2뢑s_4.��k���t�2�wTrΗ>���ǋ�f�h
�x��d��^.���K����F�C��H�����٠�?9Aݢ�]r�M	�uᲠʑ��H��9�| ĈV��A���+���V��w6���G�j�W��Ɓ�rh��ҥyZ�U���NC3h�dȭ'�.�����E��p}.�А8���e�:���3Dp>�2/E�]s��mĘ�_C���Z����!�㯍��!%��#b��ĉ�QQ���W{��"@IM�F�t]����JC�n��yW�3ב��a��I�]�ve���m�ʭ���t�Q��u�3A�Q���iس�VQ��[aˁ�r���>d�$����Vm�n�%��}�G�j�,VF��D�v���_��
Β9r��	�c>3 l���r��0WG�3GZ4Zeї��<�w���U�>g���]���"��
��F`��i�٧���p�`�����hQ��O�T�Tnj$�{����ܥ���y9!��+��ҳ��c�5f�ՂܼI�#Z�)�Dx�[D�����<�t��)��G�u4��B���r���h*�+V�eړ�U��_�4)�����؄Ę�-���D:W[kr`��n@x�S*&�Y�3�����'�� ��B����i&�t+���.2A�ND"�d�-Q]��<�Tٹ?�Lu����@���kC�+]��:����"����΋L!)&���+�2�N��\�!��_9}�ٶJԜ�ick�bV�����#	q�^�ݷ#�ݱ2nȚ��o�T�[%[�Z�<�(~pZ�zs�J*��g�������q�m�8�ߊ)�vş/���"rb�Ӓni`;��+39�|��li-c�{��.���y�d�a�q�U'�Ԋ��u7��������Gϡ�� pN��$ �qj�~ c͋λ&lD,�{bv���݇�+����c%I
�"�nWu&�\�آÀB��{�{���-��|��gH������uQ��%���b�l�P�ܜ��*��m`t)�r9S��	XQا9Z`>�.�����rּ�'�G�!g���jV(9����sd~�* �}��/=��}�!W�y�����cY)��:c��Y�t���iE"�I��C���A�)�J�M��Sl�����O�r�W.�_ �����P����k5��P<����[�#;\���u�a�zם/��"Zޥ�8�{��
b[�ww ��8[�cNo��)��l�F`����]�^+�?U�W<N�kO*mښ=�m���b�Y��t8$�7�{߁��D;���NA�dr����p�R��K��������Eޗq��֔� �r���Q�nف��cn1�qn�Y�by���~!o��d��b|%P��ݢ�u,��%3�������W�õ	���R�~]�G��,�
Ӥ�ɍ�Ima�;(׎���\jִ.C`����/���e���3/0��v �s�=�Ba�������鋘,u'��	���Y��,ۆ�����I��UKj��#�3���躰�A��@tF�:�A�0�7Y$��<����j�b� %n�	"şi7���'�NGH�&��q�A�z�uY}3<��V��۬606	���#uk�~]��}��C�"�^&��l\���sڱ�:��Q��0+������Ղ�.%��ص5�w�U8�,�ט�z֬���`Hc��UK�=$x�+��7�9'���1OI�%g��!IEZ���^���������'�ee�K���2j�C���)��'=˄�dVIN�(��q"l˨m+� :keE��"N��L�2��M�C����V:3�yRv��
ͳ�,�f��l���[R2��l��)�dh}�p�ιY�~��(m��[.s��l\[�q�ɣc�$gl�!���P��z������dp�����5xt�ɫ�}_)G�"�*^�f �2 3$��w.�wuBk�UЮ96����m�힯�I�6��n2/�t�I��4>�b���"�q��j���m�T;4ʵ�hH�0Cn1	�tˬ����ɀ����C��7J6��} �Ox�+lv
"�7�6��S<O��7��ln�i�V��\>�d��>�(�~���5\��xZw�Ƅ������]��zݙl����c�إ��Ϻ1�b?��)�!~I2���8>@��F���~���W>��aGC�RW�{��1�Mu�?&��i{@���w�r6�'�C�B��*�1EKs��Z��8x�'6�ç0��r�o�0��6�ɧ/�#v�uos��Ѡs�^����$g���@��/H"����!�ןK0}�h]�SF��9i�iP���S�-Զ�ȶ�󠂗eBQ�I���%N}R�Ku��ez�B�#�X���:���!3
I!�����>�V��Z�}Dn�)BTv��q6\z���a�;�+��q-$!~Lx�kʢ7��h������b4����E^�7���ɐ��;���)���_ �Wv��D㤃�:��U�t��6j�I���0Okԁ���l�#K���Uނ�k�;�ľL�50��4{@���A$��u�8�}�·)g�$Y�Y6���F��b���O�)�՗O��&��Ѕ-�gp/>[yD��z]�����\�CN�qC��}�a^��RXj��u��m������#�Z�_�>Yyc��F�մ]�`0��	"�������I����/��<ګPm���d18�릙��`_١�5��t���)=�Ǻ��7�q㦢�j�_n�U�'�S����m �l3�0X�T�����F�$?C���A�0|���|�N���籎�aISҚP�"fd1sK��u����'�׻p�U�&�%cV��?����.�S5��p��͓Y��w�b8�G����Ȫ�+a��j�SIz]���hf��M�b��� �[p�X�B2)��G�ː�֌�hdj�oI�2wOc�yæ\.�;�C=fpvf$�����X��l$���\])\|ɐ� �+j��������y<�Z菢�qE}޾�o��ҙ���a�~�I���?�v�8����L��?HJ�0�5R�6��b���%���s(l�g٬/��u�~Ѿ_����S�0��/�֎��}y���ކ�G��'�|V聝`wȉ�o^���W���RaYӶ�7M1{օ9#��d��7Ӱ��@!hd���)�B��|n:	⡰��#t�����?���͔C�J�.Np�9BQ��ݡ���q�:��X��=�J�	}O��Kh�:_I�Zm������r��D�F/����r����g�Wa����(�pD��Æ`PW1�4
|�|�O
?�FM̊	@���X��[���ǈ^��̴��3\ �H�{���E�.�K�G�h�v��6㚔�'��8�4�B����E���Q�]絜y� eC騤���.�!�^*�ⷵ��pQ�c8�n�q|��\&y7�H/�do�����8��.�������Yp���:�rʇ�n1I�A�I���V��o��xq9O瞅�L/ZGU-��X*��ur���TM�
�ݩ��vWRm�u~ߋ�q3�P��3���En�yv�j�sP�������k��͞� Ax����f4+��8mo�s�@]` ���0Ci��fA��a�O�O�J�>F	�3O�EC��RV��u��T�k�qs�e>fc�|ur��y(�E��0*8���5*[i���ޡ�I�J�����K�[�3����Ү'�L~J�ǚ��&������䃂��y>��W=�����WN�u�/y��]X՝ OPf��=Gx&�t ӽ� Ԥt��*T� �u��T�[PY�v�� ;���������P��vk��u��5�	�͉0��Ó�&��F$A�Ԛw��F�ؕ�L/�����c��~��= �O<�������!#�~��y�������jT.�m����J�7a��<n�u�n��|�����h�h����X5i^k ��(U�S#��{:������!Q�Ս���g�dX������6.�ο���#e`@1i1*���i�1��#��P���;��J��IsꗂR�OMC������OBpO-�.�YJ�tʲ���e#b�e�~	�O^��%������4v�q�`�z}�=5��-?��A������c���V�a��D����'�zaغg����5�"c���
��0���^(:=��j��9�^Q _�$�U$�Zk��?�	��(�66؋����6AFk݉��#В��e�x��ֹ����@����2�S���Խ�X�Y�{N��+(�8�f���ȞZt����5!jL���)���t��Q*d~[5�ི�<J��)��ÜY/���~���P�rw��	Tl����&o�u�m��%� ���d��:�]>kH����ttG�<V�e	�I(���f���� };����{w}9����r�t�?��`�>-=�]C��{�YZ�Hf��zAު��6���U�bO�Vur��oh50~���%�g���o-���p���M����Gj�CΉr�舂xQ���ʇ��fF�{��=�lR��;|J�W:4]*M��tB�E<.B���2݀��&L5H�n�^ �:�A�]{PS��/�����v)�N.)�q�Y{�����(�/�~j�_����Y�b�A5�f�צ{������o�y��8G�n[jQ�_�t`��S�K���#�ܑ�EE��MV⑒������ޜ�&��|G���~��0�����?��_D�A�w�U��4���m2�U�O�~-4V��A�'�%�.g)0&��w�gz:w&���;�<��J����0�L]"P�������58(ٳͶ~��(M��Bgr��t�y��H�.���[�hŀ� �l�f䴉(�g�U��ߓ~;�i�nB�����L���.�L��-�!���C�y�Dd�0^EG�j��"�;�`�@�@�s^!qn؉��=�L�WU��1C(to���s,BX��u��o���ˑQ~��M��w?M����!�����WCRW�DU�^�)��45)�x��u>DT��r#�j�|�#����N�b��)�ut�q�S����6�Tw�3�Py�)�9��%�6�Z�Eb\k�Ay��r��HyF���6`y��Vt�L+�?�\{�w��ݎG����^�YX��O��T��J�� �^rC��4[ڃ�������1�Ck=�'��	���vo�-8r��&�Z����j]���O�@aV�/�֏�2�Wq�蛇�t��S��܆tk�
5d��;��aF(�#3�5��ɳ��ni=�MN-���,	�O=t�h�.����?�h�$:lE��@����|�/Q59�7�^�@���u�!�lu%���_6�	"��F4(�ZƲ�e�<��A�Τ��Mp�3�IW��ܡN� ����Ia1t#�y
0��Rݞ!{ ���0f�!��8���͝m����X���jl�1đ�4Z��wr�|�l����A��K���c�zޞ�U�1��,�X����<�LӨS�Q��}�ޥg�ώ�҅csx�X���)�K��y�!�m}����5� �R�I��Xl�Ų��e[���<]����ù�4�I��?w���P��ӓ�����QC����{���L��tԲ^}ŁefLs��14�b��#k�ų��rI�� 67,�!�-C(_>�����F{��04M���q�7_{%G�f9o���c\�}��e*�ZN� L3�n�C��r�]�">}����$*��C�A]��U�,���T�������;M�v��D�͏�P_�[�i�ɔn�
�*�b�Ɉ}Ȇ�H�&_�IPV!�Z Ү﯌�;����xX~�Pa�7�C-�T�,��8Z�P;�׺Ą�ڃ}@f�Gp�w�m���u��/�E��V�����o^TEu���.��Y��a�eLF:��RS�!U���6�m���J����nP���̪�ۿ�93��F}�>≖QQ$�m�${Ž_���xg}��7���0j�<����8X#��g�׋��S>GJ"�%��0xNI�C��z����԰C�	�����f��������b��L��@P���	)ӺTu�����eC-�Z��� �YU�V�}?�Բ�H���|O�}_��oxH�� ˞[���]��s!���T�밷���9�N�_��<r���GUp�� ��w&G�*��%�㻧oJ����`k  ���'���Xd\�8�rӽ�5��It�峈:��si�%�4�o�!���o��J�B,
��j�{v!4ʧ,���\�{ÃHYK)�D��J�6)�@���hy��M��믄�w5B�-��Fɧ����!��Y���3�f܀���Ȣ��ۧu�'%�1ٴ�6�Ԁ�����?u5�;PƖ����3���~�X�S^:���uʮ_�&g@/Oa�����k��r�Fly�5�B)�U��dB4'�Ieo���h�atO�4j ���TL��\�c� k���b���9�{L�Ps`����O�I�.��c�s__�k�7�߆�p�v4��&b��֥,�}i��I�a&�����k�}��m�����
�~��"�q92�ت/�[�K�p���FӍc]~�%������%oTY���Xz�b$؁� '��*� Z�e�2p
���.D�:�QS�o*�@�6�������ƞ���R�E0�Yo����2~(n�,�l���l�O�G��,,2	ǰ#][��LV��G�ߟ}�U���d���2�@�D0��5�T�̆,M �~���!�&��q�� hk��ˠ}����Q���b��<��7�wήĂ�����|�:��O����4_ȹ�_CQu�+��}βǴ���_-�_?%��x��y�hl2��z^{�.�~��[j�Z"�ǧ��Sh"�R>?e2���+�ED����i%�I/l��Pb�ۺP�P�J(3jY6A�'Iho�y����������TPhJM�6��_Y����8�ǔ)*��p�wy�SL��?Hq<_�����%�D6���,\�D$�Vs�DZto=�V5�����+��w�T����Xa�{���!�Q�%�z��R��(�4Д���>Q.�7�Y(G��v<6�����-'Qq���h����	U�+:�Q��F����6K"��0�������h���7mv��������1���� ���@-|��Gqg'�M���E�w�m��ijx?�9�ӂN3��?���#�����$����.�s^��V#)3:s��	��?Q��|��
WM.Ԅ`�X��� ��٨������y���N���
�m����3g�+��*JT@��5��X"�Rn��Q�����Va]C)a�B���=�����֒�WFGUG؉�����(����gk�V��xb��W�;���Y���������j�rR!n��xl8ᠯp�y�E�j\� ��Y��3X��/t�y���!�{���hV�|ssx������N�znF$���RS$�@T�/�T��R�=? �<~�;�\��w��>'d�9��fIs����0=1��$K��T��翷���F;�-�.#G Z5E��s�H���{VN������qV�Jys��8$d��loj��"><�7Ӡ�Z�s9�Wu�dl61��sd��\��G��F,�)}i
���]�Z�8?r:�͗6��ν�;���{�j�tw�"�+q��װ�
���2�)�ΥC"�]ǔ� \@�i�J��1š]��_E�Z@�d�>�B$�|�I�BWƤ݅���H$4Y%�ߢ%5BIa�J�JjNgv���'N�����F��{� �����sv����uYgN�ؤ���+�`��2�$﫻m-s��@���ۿ{�&���#�M��V�F�g� ��(m�y%ܬc��z敉�~Bǲ��E�� ~p�� c��
\H��� B���e9��(,)�8L�?2袛d\&#���~iO��$��mф��4�g���z�Fc�a�>�xf�1F�8
./I����)U~󷻜Ѓ�'�8n1�Ж]i�{BFF�(Œ��2
�k�Nvɶ�pV��%�t�D���>bJy�ؑ�?	ս��*���$�0�M?���]�!`!��o�t��56���M�{��T��\�6����0\�g���)�τ� ,3P�,GEl12QR�\ʯ�5�s-�l��T,i�~�蒩��)�f��y�8��Hu���~�5u��oU���A����Uk���qk2rI�~�������Y�PG��"ŗ�z}g~f��[��L��`�q��9z�S1�����b����c��!X���j�W/�h��P:q.P|���w�������`n�"�G����A��x�`:\��nQd��+�x\���4�[�4�`��ay`�1������fO�{�@�ͮ�o�_��]�� ��WR���G��BY/d-�� ��.��AC�3��3=�������g�E&�+��2���|��!�t����j��G`�2��1~�����m��>�$�t�_�1r9$�����k��r.���>�YK� �)��[6�J��Pf��?u�:%������$\�A�<�5�pcJjz�J��^w�vTuQR`F��M��c����Ͷ���KC��E�m*~WWd'����w�re�]cP�H��%M>cɱ����*��}�b-�,V��-��j�A�����gW�SY���>� }�sG���R;��j���$C��@LU'==��^�E:�>n31:�!2���=8���?��]_�N�������	� ������bʯ�P�0��_�O��i�\�*�P=��J"|d��@ŭ��~4���IA�v!x2�\߷�'ĕf�tL�k(��W�5MJ�ƀ��_��A2Q��#�	$?e/0�����j�뛾{,Tg���-�!���ZQ���6m�[+����Q��1�3���ؑ�ak��7\vd�l`��=�]���+���\q���VJ��B4 N�b.0�bc��޶x��n<�6=uN��pj\��eo�i�	i���&���]�e�_/Ɯ�ȁV� ;sz��9���7�ᮺ�+���רw�oͤD�It_+8��ɼe�۾(E�0���Iz�����ٓ��Z�[���1�f}d� �&'ɪE��<B?�Q���e��^t$�ƭO��#�b�u��O��-h��ވ��RC]ܙ7�䴤^$P�ս�>��ì��S��"��I���t���嶿��3��NI�fj�*��&ss*y�$~ �Ϙa!	��=�H�d��xwⳐ4�sSW���,Μ{��Q���:��_��z"���"ݷ'�����$�Dkr��OR�����ʸL(��%���@��D�/�87Ci �&��bN�hJ@�K�����r����`PD؁Dd�Y L0q$Ih,Ͻ��i��=�k�wq���Q2����V/W�X��2���9<[ )�C��ޠ �_�:Sw�K��f���Y��=`���a���"�1��ަ��?W_�l�y�����t�^���B|�(�+�vB�C����j�q�#(Q#|��Zo�H�.P��yV/����]L�C�-�9_�����"�C{�,OyMg{+�����d�Y�6i��r'Σ��>�.5�!g_>!Au�i� �*��O��sƁȧz��m�m���+�NH���=X�2�(��8�����z~���Wy�G�������Jg:֕,��y�Y���54ERt��Ry�6�=#��3�h:�t؉{�:H�=�8:�2�Háͼ��r^�#�h�����S��9B��i�yhB)s�p���".FM�Nc�Yh/e��^=�,(��-�3�(.�ޖ6����y:�J�z"#'_���]I��>gT����GT��V�L0
��`��;�h�=��F����0�����T�̹N��,�)S�1���@�͟��~/>} j����J�>W)�(�mA��h�<͑�j�~TwrۚYg3z\ra>�Q�V�����;n\5v@�;Rǹ�a�	Y����'%)��[(PU��Ih��&�bnWʾ/�V��*�����M��&�:;���m�[�<E����BR�}���|��Z�Ȇ9 3���#5��ޫ���D�ٵ�;[P#��m&+?��`B��P�D��X����F�A���ͺ٭��WG9X/h&�\qI�Ӈ�ǠSʳH�/����U:)B����<8B�OtZa�����M{TzgC�,�~�G�^�?����ce��
87����O�tEO`��;
�팕�W�펢�
��Y������\�%}�CPR���7�7ӊ-]g���'�CP&/%ъ]��#�|*5�Ʉ�҅���Qpռ�A�x��
�0W��������`��P��@sf.�����磭��z�]Ю8ѓ���|�����GשY��Z�,���B�{���@�ۏ>t3t�P����~�@Uve��tw{Xh��v��"�&��\Mr��;6�s�7_�9���^i&��k�#L�0��C"m5�]{�^���
uU
PG��4�8`�{�G����	[�� �d�1)��߹�?��F`��V��9@����\:|\��U2"y�q:0�@`��±��O�i��	ׅ_�S�z�������\T��?���j��������S�GX`��H-HnOh����V�
�|��-��	�-ּ>��ZUr8�`?����TK��ṋ2H8W����WȆ�Dd\�M�O ��gJ���b�\�|�˛g�y�l��䙺��9�ٞ���,o�M�WS��7n9H�'M�1R���ᶗCO�rE�L�OG��D#^m?��W�BO�5�?4\����R�NXN�x�,�>�E L�>�EWv1��׆�O��J[�I7KU��q�h�Ϯ;[y��>�O�N�n��z߄ӫ���=�}4�y�p�����}�}�����%k(4=�hG%�P����Q���)���fl�O����;�����[���~�U��|��nۄ0/=vB6���݃��>��{j�M"c���~��:N�.s��%�k�!48��Wk7��ᡤa�89�-xՎ����᮷�T���\�O����5t|�E�gR0F�r��|��r����k�ABkUC�j�U�悌3l@O��<�,oL%�>����AAI��YB`Wy��?sXc��c�,�0Ѱ��!Nq\k�/��،���1j�P��>��8˕r�ZX  vK��I�rW��h��2M��.�)4��P��.�qS�(nH}[��NJ��Ԯ��S�O&��R˪����Eæ�x��h�ꍪh�Q!�n�����m�����D�8�/����Gܘ,^�|��.���.�.e�C�d�����ӗ�:=O4<i�����p4Q|w4�P�s�<����DC��$bp�zѼ5���LU�F�j��p�E��a��<��CL��=ax�q 1�#�]2�F�3_'�Tڲ�I�LlJ�7~"�0���U�9�S`��gŶ=��8�� �0("�,~��(�1}�|�����O����"�T�B�n�����8���M�ިv��Q\��PH�wm���4d�)wW@8�̨M�,ٰ�kpN�aܫVA)|�7��x����w���:4��Lo�`��K>��[�@���-���9����O/iX��":�+.&>�jkw"�k��f��X�Ӵ2�R�i�tP��!)S�\)�م�	l �[�IV�+�Ѫ=�v�* �������<[��L��mJ�_#�������ZQÂ�ߏ�p�ȑ�1J4&�!�Q��XF�&�s�$8�	�06!?=�qΝeCeB��\�Gy���Z�XIkf��/�"ܖ�+ņʲ&\�tg��p�aҦ���N��-����e�o�}vM�LaNUf�;#��訍�?��@�b���z���y� R�Νv���[�5��w��F,kqq�e|s-����#��&b�S63Ki/\p�����G��;[P�
��D��/F������;ͬ(ɖ�S��*��-��h���B����@Ik��j�ii:<q��F�r-�\����boWlg�����Ҭ����S��Bj���|���Ȧ��n2���X�R� ���aR|(��@�̏�Ӆ2E>�x]�HD�5%P'�&
6�l���Գ�d�.f��d�JD��H�^���60l.���V�o?Q�'�rjt��x��w��i��"�����m����~�U�B&wQ �4�	�����.$Q�~ڋԜ�qK>Q��D�l-%w���$���z���j�ݬ���ф|>�)_�����d��a��K���9�h8���_�Q��|Aˑ ��&��5�kv|'X��kf���"�£�^i7����[�
^
�t�_�e��jcR�%��]*m�#����@ɸi��X�j���_k6�4n!�j-:L4��=^[{��a?a��{�:ry�=��ю�j�_��6���`v�yWW�p�U�}H�O��Iq��0�&�n/2��F�Ә�+����",9AL0�d�;���g��!��[b��*�D"�K����9d8�	E���M>0t^��tI�G��?�����!��^?c፴;���J�[_�
��;;�w���h������s-Hž��b�0=�\���u�qz��� Y��׿��{�@���dp��#���i�?S�l�#�C���Ȼ� �v;RR��L��m���(�CgF���e���g��\�V�l�'��q3<�Ȃ¶\��ϗ��n\YR+�;S��.�G8F�Y?��xTB�[|2ji^z\�� ��ۋQ*�����P��5i��V��'�KQm7_�B|Y�>���y��2�.�jIm��>{Q8��x��|�����x�G��Aogz�^BgC�n:
�������tĂ�I0�@Ơ<E�
�*8fK�iA��}�4�Ƶ�M+�T�ԃ������t��TQ�;�k�D�-�˕(A�'��7��C�UaR[+*�g;&����|i���t%)_�p��ҧ~R��,��;�1=v��R��W�k�~�N��WHp��V�Y'�.�̢�_*+������|쀗
�y��x�C~��;{�گ}V�%��s���
b��:^7�֎� ʠNh�i�c���i3�[b8��t�b˻��x#'0� /?��� ��ú��.��[U�5=�o�}��������$_��37��9 0Tr;F��)Ќ�$��`<�Q��@�W��=��\u�Zj���;����>�Ã�f�s)�{ZC�A�����P���5i��@��5@���[�~�����Cf	�F� �}c���t[���U(c=E��su`5]�0���1��f,�IίDB�6�tc��<��=�[)cq�3[T !%Xe!�U�J�����N_�z�I�S���xU�������
Ć0�J���yή�r���r>�GI,{?	���*������U�x�S�%8�0b"�����g�ז��|w(b&�%V'�����U���`�Am��N��_ |��𣮝��{�!�2J����7�}6��c��Rtzf�j�p�2�.*$�sU΋(xo����a�{2\7'v S���|�c�̡���xP�� �8ߦч�@ �rUϝ-%�T�N���=��R	o1�f�n8�DJz���sV"j(� ��
�5�р	��,����p�pG%N��;.~�X۫��H��jr¡ۘȵ	QZ��N(Y��o�g�ra]��(;�O�K\��(6-&��D�4��oO�B�z ��oW}!F~G�v�	ʱ�v,�k!�/�:��s�ˇ4�4�dq��U �+���� XG��3�j�K���0�2;[��������W�%�A����m�>����=ĉ���m���터-n��0��" 4�ɹ�n�:Z-ѨaL_���Q�	���� Q������1B�����l��_�w�d>�w��n�(>=�ε-b�e6���K�j(7خKyq�रc�.R�Q+ �̯�!�:�%��$	4Gu+`�Z_��uB���g�7�R�l/�c���cudM�A) ��:�h� �7Sa�6֝ ��C��/T��W݇��M��C��C���;�+;�lz�ܣ�,�eM��!��)�R�/���y��/1�9���Q�|G���|�v��׶�i��
��)c��C`��8���g�#)1�ڢ%�-�Zb'h}MJ\ld�thA���FV9�.K�@��(}��J����W���0��,t2,�S�ߩ~�y���{�Hʷ���enk$c�G5xZ:��Z�w�bH ��K�'�������e)�Hz��[!��h�:D�=�J+ơ��4�>!_�눿E���H����<Q��� ��}�&0��D�TOa:���)0h5J��9��:��"�A����=C�u�Ws`r���tC+���F��쏲�.�0u/T�@��8��̮�����x�$��5�϶;��}�/�줳e�{�ޡశ��omH�f�[�
���\�8�� FXI~8�Y�{V_4��-6�D���qd�J�Qi�u�=��i�sK��Զ�Ga�]d��"����d7���T��@%�{P�xW�حxͧ���SB�&ɭ�#���,�/�z�(��$e��B��ȿ�y�V��R�B�	�C���*���cJ���AG"�.o[��������H�h�T�ې�˚o�58����ǉ+2�PC���\�R�0vk��e� zǬ5v�����@�~wD"�m�9���M�U�8~����*X	���18������G���dz�(����a����D��2�xo�M�`����&MY�}۽�N�dN�o0�Yp���k���O��l�"a"sy{?p�M��\��;�Ҵ�*a#��w��K�V3!���G��'��
��i1��k�t�t)ө�q�B�}˓�|���Y>�ͻ�8cլH���ux<�tCY7j���,b��34-��~l�����a8�zO�XJ�y�E�I�����$��8aK�t���Dp5�Ür��`_w�t��nn�h��O�O�Z�ԁ�˷�m:d�hv��Y����h��A��az��M�-�hoPw�|��2:<�38�A�7��q��TNa�J���k�&6�/�W���RÒ��D�hQ�o ns��c4q�:�3�,���tUR�7ě���ߐ����rT��^\a�q���� ϋ�@΢���t���M�|������7�� c��fMf�G��������uW�3z�a!�$�ՉD_��U-~7�����5�258ڈ��J}��՘(�0 
��y^0�f~������-���Zռ��]��)�$�d���Hb��(��3\Pwx|��m�	Yr���lₙ�Um�\��A{�7�|�AhD,X:{h-���މ���<�RR2�j��|_��֋��ܖ|�לw�+c�2����F��O�&3��-�f��G���]!=�(��ۘ	��+~��0�A�/fb�ݚHW�l����I�?��l7��+W��
��b���X�������r㟏�y]�V��V����Uɾ#"�%zn���&��h���=v��$�_}8��j=.A���|����:�=�*�]�nQ��Y~��v��a�Y��U�4�X&�~�T�y7Λ[:?O����ǈ��hZ�Bx#�&�kb@fғ%[��qr�y���g*I�� J|���;��P��i-P�uE*7�FkĐ���35�HR�Cm;�����;�yl}�c��Qn9�-{��Nf��徵};�x�~�h��P�R�����_sU�aC8.0/���x�T�g*o��=bL	�~�^�F|)V:C�B6��D8!Mի�
ׄT[��k�;��"�C��>A'v�.Q�]��2���^��������qi��1�'��^��Z6��'#�B���fk���KT������A�MX�?�o;����g�Ω�S�ހ�Nh�Ӵ��eN$�|Y��:&�0������R��w�g��*��_g��WÎ���A��eM�ϓ7ŕI^����$�a�-���wu�0,4V�=��A)���wT�n>μOjG�D�J�BH��IwC+�w��)Ֆ��cC��n���G�NqfT�HXZ!�-�5t�,�W3���A����V�����[���g��@f�d��Z� �h��5�&�Be�`ʼ�HSZ��t2<��Õ��Y&��R݄�T 7&���M�=k���'��1�Ɗ�"p��q8�^�hS!����L��ϦI���s%��"Y5z�었�F��Lϐ�dnζĐt	�/T)��������f���#����f�\'J�50`�:���"����M����h�:ێ���?�J�����жu@>�l����d�R�V�ch1�n�PEӜo�����0��Vn[PvKfT �,#j����`�}}ƀJޮ�{n��x���j�20���o����;�����'��{��W��@�,�Fp$��b�.�_��U������vi�Y��Bg�n/^��u	a��@�T��x����Z�0u.P=��}�[/7Α�#����\	A�����8~%�����m_��ڶ`��ql;��	�v�3ZS�0B�T�D����g�[����\gdP��a`�\�����h��RZ����!�����v%�MF����{d�/�e&>���ɩDK�iX"�T�[n��1�i؆ȷ�tnzs�pK���ǰUߕ#� 񮦐:ChX(ҁ1�S����Xw�N�3�S�'����P#��J�?)�b�fo�m���K�NX��il���E�X?�
��:1L�Gω�1�����ܳ^������.4��@Me_����V��3��&���j��kc�8$�������,�dN�RQi��U�oJ�EFgA9WvI����bP��5�K&kI�{{�2v��P�W4k�'���������ޡ�KUfFԻ�`�'� X����3_����u�e R�3r3�]7 vX�����!�����BQ�)r|�&�������2.�7�H��׈܊}kE3mխx\M�>������j3p�q����W��m�f��Ҫu���.��3tރL4(IY�D(*B�iv�s&M�!�����K����J�,������j���8^"��FǾ��W�ʱçi(O�ac4j�9�`��r�ޯ��\�@ψ�U�"�=|���Y�y���U���NU&Q�qQ7�7S=���]�~iUtsu@��6P3���F��G����+#�p����9Vh��\8��r��ACa��M��h`*���cZ�o���XY�8�,��Wj�#_���A�_�X�,�(����9jVT�ODf?0�ʼX�&\�V<����+����5��[�[x9Q�f��U�T���
/Y�3z�-R"�
6y�މ���rP6,o)��TI'^��'^�cc�2p-��N�����h�y����+)|���}���B2@���Z��ոb��b}5�SCu�?��&�>��7/Q��y�t}Q�6��_�����M��D��pV��S&z*��MI�zj�K�H���^m�CaÃs #�f,>�䝰�F�P��Q�6����^�����$���3�=��Rf@&�n˶�׍�"La��FNg:Oz/zY�g	�Dq�g��u��(���>��,���Y����:�չ�������`}Z�����-�������7�'`�����>[ RQ�,�L�Df���/\�d�<m����]xD��qN@�h(�:��<��?hf�>��l`-�<����ʜY���&�e\]�����
�(�Q������r�O��� ~� :1,�e�}3B�fb�_G����&��5K��q���X!<���W�
��D~��Q��4O������΄龋�o��A%"TjL��W41�(G|�^�5ږ`�w#٣m����/&�������Z�^Vfo�j�\�S4���5a�����G��=t"�+�fΥ;��^�[�S�LEp���^��vc���U����<�R-�n��J���1$$�F�!��=�8R�5���@]��<($����L2$�� J�6o�;�(WN�Ϸ��w5�V�΄�(X�E�HZz�x|�,�*_&�9�u�����r�+?�Y�U̯X���~�)]���=G�B�w ���nV��l���G��ك_E0)M5��QaF�/1�|���j�8(s�	F��i_�!��،���˗6G�b!�|;���y$<,s����/��U�p�:�ݦ��ڬ)b�VW�aB�X/� �+}
�.�c�z\�A9B��R�(�����r��bs^�1��r��	�H�њ�Bb=��/��T���  |(}������������h/�; p;�ït�E�5t�i��wh��뫐�E�a��E�f�f��`�q^6[���#���_)����j%p�wМ��՚��Np�u�f�<Xc�C����PY���3?I��4��?��Os�̻9�I��y��}"D���[fm�1{}�907c�'��|v����lτ��3���E`�'��$��	!%L�ݝ~�[�#�N���QWe�� A^M�9H�u�4�t~'�wWO�&�T�[z���������\�ž�R��s{E���q�;����MP�RHu;��u���?iiĻ�) ���xxǕ���W(B��7��+���N�娳�	�Bw�io�d�pG����
Ɂm��S�?��6J�#�����5@u5� y�<�:i"E	�#�2qi

eG�\.��+��ԉ��-Y�f���&�</�}�a�\�>{������)D/���i�~��k���|���豗�P�i�]���5�`�f�ʒpn,%G_B0�5�n���Y���ړ:t�a#F�?��tI�����|��O�:�([��RS���2��Vh���f����kPӂ��P�)1u��3�Qǐqda"�����X�*�	{X���+>����R�c�2z���vҭEr�s������(�ِ�"~":��Mf��e����������秸�YH���@�zũ�"k"�`�M�re1�{?������Y:�ܨ��̎�q��!���i�<�,�4�G{bR��g�,^!a6�9K]Ŏb
����@�;�|䊾�����p2_	=�+ۘZ&SA�-��e�Ig�$��"�
OIh�Z��*jJ��!��zZ����9�'�$]�9�q��/�c���,C����<�7&���K�ĸi��"��<Z3:d��ږLO�>^K���}g�XN�R�qj��ɺ}:���U�")�e �oQ�h���Ma��1�T��j�HG�Q5H�F�/ټD���s3�j+7&�~B�2��X��c�hE|CA��d�J��猰�׈+WBÛԖ#���J|\]%�]���@�A�Y:C��eA�*K���W�al�R�h��>��6Ŏ�xu��V�[V��c|ӫ}��#'$����[R�	�2��߰��\z��[z?�1�q�T���Ziw �ᖾ�i��e���΂�-gz���7���I�c����x�:���1��c!Y��o���*a����I�6q�T����\k#��k
�:��n��s`v"�=��Ș�Md ��jU�z�e_�B#3x;"�����8?�R���F�b���B�;��*p<m�ʄ� ��v�A�����O� c�ǳW�;����2߹8Ҵ���F�G���Qi�N��:�u��A���b#�/�A*<sq�[g|��P�������l����4�%�aG����"�`�,A٩֑���G�_q���ݨL����(���"G/k�cu�1�
���:�a�݈��x�J�@��fBl��EA�}��ޢ���������3$Af��u���-�ٚB�BT�VW�Y(wb�G�ZR�E��v"?p(?
�ۙ��@��kF��1�Q/Ќ�����5m'nQZY'�s"W�B}Rג����K=RÖn���I���>N�����^��a��ѓ��<AAEd�5D���1_���j@�0�n�	Ly�F�o ����^�k?��,�M(q����f���{#<,D��Ӟ�mkZȶ.?h�
�&`�� q����$�d���L�3�%��j76��hNJȞ��\�2D?:=�B'�x�J�*��Qٽ�5� ,��Z�Y}��+�*�0ރ�R��g@�������(��LĦ~�!��PX&z���<��
��y�� �&J�3��g������J��p�lh�.E�������ۏ�I�����MZ;T#=�	����������n����׮��mYn�B��LT��^hC��Y�6�r���$�J���B�`�L�n�v�O'��D�E��֧��O�lJ��:c���{f`Vߣm��S�o�&ت�s��-����3gS������	i�B�ߦ�yi���PP�!e�*�(ƚ�L�Q�!�\��e�Qƥ4�b�f�s�aP�iB�����O���SC� �Ka�,�9)�0�-8��0�/�����&�&�N^K�h~��KZ�w̉/�/c���ֿ�?�����m���]Ad�q�w3:V�a��Rt�Vl�-Q	'�j1�@a^��'�e��p��[*�0���ť)�,H�@Q�a�c�?O� ����zƊ>�G4�i��D�J'��ƁF-#�*��������
���C�u{\:"�����h҆�Xb����Lp�@r�=��jY��+�Ռ�.3�$-bV����m% i"�?K?��WP�5�p�Au*ω"�J������U�wun���		D���{O��洠8��eF��NK A�G�+��r�W{��"
��U&�!���F���AhV���Χa9,VJ-3�����U�F����\8Į�����T�o�lgiy��_$�V�ʕ�tc��c`$��C[C1S�#���bTip��C��"P:���t]�[(�{5{Q1���5��,���s�Su@$� Ra2�i��0��WT�G)f=��	�ߡs_�dKQ�Ə��QD-��{���o�5�M�A�-��D;������n��Y�tӭ��Ni�ı���7�d���5���(^^��2x%�yl}���7�?Fh���3�8 A��#��o��� ����4Y�o@�.�t�6Cg��֐���70<��1߷���o��!�`*�f��M#��b4�o���0=5[���O,��g���r
�A긣�0tJcʚr�[�60V6ُy �t�jJ��M�#Z��M���h�2m�e���+C{敾��j���hF���~�O���ͼRl��Tpb��x
^��p��N�TnT������i�c��Y�,؃���o�˦��A뒄�_%���P�	��)�Dm+U����VP�?��P-�����G�b�h?���?����c�Y�̳R\e���;Q���0�ƚ@z���5s�#0;E��h�3�1��G���`��J(o��:@ep�������!+���4�XQ�g ��ȕ�j,��P� ��*ze�kF�҃Ì�}QEOb+�H%��5A}0nu\�Wq��>������j~,��!od0�2i�{0(j��7�/��g�F�=n��M(La_�W��(�4�^�u�������!y�v�*�Ż�t+�WC*/�x��D��mƹҎy� ����rv�(P�Xl3�nK�ś��:/O���� ˑ(k�7ѬD��Hw��G�Q��5�E��r0�h�dh�'a� ;ȳ��A1���_�P�$Zs�%]8�&�'�q��aR���M�wM�3ɥ��G��`�����[J
�|���N����#��:ޓ[đp�Z��(�)Ԃg��fUh���#�����^]dNA)/w��g!1q�/�no�`V�W���\��I��l��K v���b��@��W��v�o�б��=X�n���Y���v��8�U��+���I��;w�p�E�1�:�ٹS���(c�O9���@�/`mul��D�=�JO�dF C�(�}�����w̑�ϛ��F%G�
-�UK%����eJ"������0�l�S:���E�\�������K����_as�ծP�0*�刾��(�^A�N�t��j$g�9�[���y�&F��j�!��[Y!T��25��6��k�m�|���t!.\��j��'I{B�$�-9.M�'�_ʘ����nC�Z�"�0r�Pg.�1�i�~W=��;鵝�p�����z�D\ݐ��=nB�e�ؘdԿ>Ț{������S��j�a�� �6����CF�,��=�Z����C��G0ʩ#�"'�~��B�n�P��n�2�miy�<G,�b��X���7�C�V�ZF��U�o��a�F�~��G+��Y�+�` |xH���)_�O�6)WC�ʕ:y�Ϗ��٨�K�޽H0���^��T)��_�<n|���I�ȼ>!����C�p_]���	ܪ:f'��MZ����`��g�ĦEO�8���Ϭ�K�^��t��#���O)b��%�
�pa���%���kAA�/���]}V�Ň0�[Z��N�}M�m(�%�L I����Bc=q�=�j�l��Ym�̜)�x.��kHg#z��0�h3'���g�V�	 T*�����uP���Ç��e�y!����) �$(��T��h�7Sa��xM��(
��"� �S���&��w�<{g5ir+z>Y�,/���쁽4'�> �>��Fң���<�|����2W΂��/y~0�߄����r����ᰁ�� ��-�'��JrS:�pɬ�6&3L�������Pj-pע�z��Q�*�b٪D��1>#X����2jQ��S��}v.�g;O�M�H��0	'O/�*J)�X��[0��y����Hr�Z`�Mp��᩼����"!�iD.KfD�W� �R�3 ���:�����ߦP�Ї���Wgq�ԞOVu��L�/|��: *�/�t2]й�)�xU���WrE7�� s���@��%~(��p��{öG�����i� ����H���c���rNq�y����o�QP��s��FNc��kC�ENد4��H[����f�6Tȗ+���!�R�f`jh���h��{PA
uu�x|$��
�F�{�o���cK3Z��1�H���<�h6n0�n=W�.MZ�@�/�05#};b�c!$�UɈu$!jxnWǓ+�C�	�i��>|T��e� �;*(�qy+i�R�(�e`�A��"�4p��)"�|����=�隠A��>��8�s�J@�B���q��u����!����ȟvKm6gyb�2�F`n�z�=$L�B����q��T,2o��W5�����KS�S.�Cs�xf-�ED���}Pv���첈krnS�v�����G�L
*'S����.0��$��⒂Ez=lF��X�$̘���'����g�f�)��O�����W�5�4X�ߜ�UT(���]:��X��C�ނ��[]��� D���C�1t~�@y� tַWF%�}=�٘�w��S��?�!niM�"`d�}��&J �%��*S�n�F�U��v*t	?]�Xy<`#�XQI��||�KYx�c1 �|K2P!!�	BW��h�2�����C$�����L�[`�{�U�p����~	��/-�dG1�^(K�k!,wa�d��%���p��!������kԠ��yV~�239�h?	Oe@�t{�dq���!_֛��B��ҿ�iy8eP�Fd~��mk��U]Mz��|�KR�zM�}��V'�i�TZcl�D"�X��V( �QTr�P�o>��th���"�|3�&A�f棚[���i�|n�YP�Ml7��]D�V�۳�ԙ��	��5H����Q�O��U$��f&�g�;�l�����~�����v4S4�f�}y�z���r`���-i�H���q��cP�H�����M|}�������>� 5˱�e��&���=8�����2�VbȁqbhA��ԫ��<��r���D��|�S]v��e�؇S��M��ڰ�U����,9&"�I�<�?Q5��rz���6����)��{)C4#�;��0�L�}�4;����D�iq� ��Kȶ	 ۋ�ƍ�EW=�k0㽵v�� 8FG~܈\Ij�1Թ%,�������4w�~ͽb�a�ڨ�7��~=��Jӕ�����,���!�`+g��E'��Z�S�9p������̑��_��~4��!���^��|\lPW�$��(4�<Z/��W�(��lJ����2�	ρ�+�֮��s�P�v�+JTی�����Y|X���^Gc�t^�&����6�0
���՚0d���4=�P�j�y��pZK��n�Z���k�LKn�K�+��]p����A H/!�J�y���KKP9�-L5������ ��#q����p�r5T����QjEyoq,.�UK)�]�k}�l�s	-�����?M�h��d���B���MR�FB������<Cc������M(U�4�%+۸V˯Q_3(Ϸ��Maq���T�ѐ�s}�8�B%�i��z���,�(�)do�ق��G!8k���>]�=t�ٚn��NyCȄ��R�i!4�ޒ�[��Iz�F��.���sdYQ��	B���[�`m�@U8B��M�~�s�e=��	�)���5[i�G��������e�@���S��a��n�3EX 5�!~�!-(=��-J|�#T��g��:�DY�ɕ6�V�7@۸���;�|E>-���N|�٭�T9��H��.�����@�
|E�T
�PM�����6,ЛK!�E����joh_���qe�~Vc�9����ΎF�w �w�N����O�V:^���8��3��\@{G���>%	�$J��/�|ī2C�b����WzM��4��0��d}�:V��Ð�K粟�q�˜�x%��ĕp\�~��v,��1ð�]�"WVlS��:�"M�}�^d�������I�UJ��V[k��?�UN�0=z~Gܬ�����Z���S̃�F(g_�C����~���7�.|1h���D�� �oQ�ށ,T>R�FH�����Lzא��X(��x��Ic��5�S<�ӊ���X?����B�f=J�� �J���S��2n��ۜ͝�"t���6Tvn�G뼔�%ݍ�^]�$1ye/c��`����u�1�u��c�?�'�G�E���/*2gEZ��m����f�lޛ�
���I3��(�9���C���OG�!B?q�>����o���q 
����Q�{o!���+���}�*C>{}�hM��Ra5���j�>�H6��Tk�+´����P~��Qu�tk�o�#HhJ�0�f�a�"�u�w'�	g��w$���#�]���XG���@�]Y:#�n�G!�$p$WO�%V��'�7*]��y�\��V?�OMZZ�c'��#��p�y��ٹ�GGBfC�����0r��p�N��V�-u�O@"/�J��po�����㥯�8%A�0`&v�uϕ���2zp!��F���'�?P3ta@�Ŷ�uQ���h�e��������c�"����0*A��ng��¨�}����g#�����B�Z�+��\Ǩ�@2���[�>�[	:q��I���X��.��3��7��cq�+Q^t#��y�<n�U�1p�ߔuL�1��rfG�D&���5t���בȭ�m���YU*���~�F�2瀓VE�Q�,4!�lHE%��Wh���>*j?l�8��&�	�F��{�F�m����_��"�&�(6��/� W��ՠ����"���� ���d��O�a�l�/�4��!L��C1G!����S����4G"(�m陿���
��Y@��c�§8+�v@�	���,�8 ��A���Df�X�a}�<W�̀�W���a�F?}m7@��KK�-/����MAɣ�#���r^?�\��1�2�����`p�v��S���]�z��&�F��+YĚ��ѠT�"��!�D\�w�Mz��x��k]�u3��.���*�?`.���+��f�D_J�o�7r��$��p�;��w�sҪ�ʥ�\�Er y�d$�%g�c!�΂3��1��D}P��4M�H��OTG�&C�� aM��/(�<�Ƿ=����K�Q��[F���>��m��ީ����eJT��b) �x����+�9�ֻ,�!^,W9[v ���c-�� fh��gP�ǯܤ��o+;?�Ý�����s:NaHzܰ~zb"��F���d��%��&�-(qDSW��BM�����"��nPfa�k��(|u	����L��99��A�!����<d�^��\:Hz(�C�~��N/˞�{��H�m�	4���,�8�J�
v`��T�����_I��r�r/x�������Q
:���;�4����@jb����PE�H�'����Y%�Fm��)5"{?�����sO��1\:��$��ުNq�+}0绱Bf`+���<
�d��5�҇�
����	=�S?����x���k�N^�EW�,Т3��*B�����[K�_�Y\uhXM�
���w��7`36T�L��9y���4�.�C�j��դR`G-$��XmC�����G)ݢ�\���ҏ�,"�lU�|��*R�t0G\�m_��s�D�^Y�6j�P�e����IޥC����,2�uЂ��me�����YT�7\%;`��;l#v3�t˴+�kS`ep�N�s�4E�����E�'��@C�����ig�2+ �:k������R_u �#'�\Q��s$G���#recv
�1?S3.i�z��ۜ�V���t�#��B7\/��[�	����#9>w�֚̀C��&�.��+��'��a�$e�+Y5����W񿿩{"ȏ'��g��ۨ��͋@�v�uf�Hi]�љf�֙��<�J�p�.m���d�� �.�Քw<��hѐ0�Wk��{t�ĿDa�\�̷�ó��7���B��-t� ���y����c��$*�B���Rv	�׀���0��g7��u��
-�n��邏2Z+����(2%�T��2��Z(u���Q�[;0�hu}�a�T��h����)�ƕ; B�&��S���E���9u����5���P���xB�@"�����+e�4�=ݢƁj;Ƥ���X��)t$���'�ŀ}E;0�v��`�'<�G�ҋ��+L?5K��@�nr�V�.-�v�+SB�`�ʳc�3����B�E��S�;� �L�86fi�~��ߟ�r4yM�N���{ٕG��p[�q�DmFF��;�en�͌��)pNx�˚g`���BkZ|-}Y��C���z%`)ě��ͮ�z+4��[U�~~���m�Q� ���ST�z���K�cf��@7�B�����W�����D�Ru��������9�zԣ$�G� Jj��(,m��XT|��n��M�3A���(���'G�BCG����Ы���ݬ�Y�'�zt���B�8�OQ����n�#(�<����w���.<�E����Q�����_��l�zPe�AH��e�(��ɞǚ�Cr�7��G�qRY���.�_)7���k�톄-=���wW�m�7��
i�ł�,jj����K: ¸�cF�f*L�� �Uq�����v�[ѳ&.>��ѤX>�0.�2�m�c�A��%t�2�(6���%�U?}+�7��W�B�ݧ��E�h 0�TEi�/�5��y΀=ݲE������܅3�� ы�+��G�����{l�܍6��/��XE! �����ṇ�cX���[[2�D)kn�^�	���_�
 H����ID��p\���H�����0�!��^������T�)����j�루	�nOu4ƽG�Ca"8�Pq�Oe/<t��c*��T��ȀO����f���6z>����3�� ت�b�a�q��$&�uǾ֧<xB�KX���ե{N 7
:�V��j�	��]�Pv��Q�q}0�8�a�32hN.�C/�R�M=v�Zuq�G_ya|�)aO�,�K�S��{�"4 �W�S?<��5�b�]���d��@o�b�,U��.��u����J	呩3bm���FƩ=�����	�&3 �����y��8�G��w��m�)/�0'����Ӫ�/N�Yꢠ������]�w!8aT��Y�w���k��"]%wꧣЮ@��K��N"�/t� �58�@J�\�8�	�Q4ˑ����G��W�8#J6�??<�0]���w/�"n����w�ո�צ��I��f3G{�c\��Y?�?W.�6�co�!V"q\�e;ݔ/�f=�~����O���u�6q���@�\�W5H����� F����+$�:��-�*]��	QJ��}�s���'�jjcn@)���	+�uR�|�xg�J�ͼnJ�Z��)�Ӳ��\ d�t�:�
��[u�����7������
����a�
�TM#� ��P��E]yQ�$�Ȕ��W�����n)�a��j_}����|3���e'�������q_a���Ñ�}&I��l�I\T��cV�)½�9��<���B�����݉�4,@Do�S��	�Օ�L <�����Q���QrC�䐰�ja��p,>��c%z�Ge��gYa!7�m��� ��e�~��I��Zu=<I����R58�@ri�>�s�֌�
P���Q1M�q5O�������bͻ�F�o�	[�N�Rߍ���HF
M6������Z[�y9���"�Є�g8�篗�aRc���Ƃ~�t �II�)��,�q��-'���!8����Hy��zR��3hW���	���,���J-���*g�T����S��OV����Ȱ�5�b?��䋡jE��b���g �]AJr��e5�M_�
_��E�U�	¥��VrA��v�KǟȊZ��^0ӿ�·0-�������U »U�
��%/�L��o��쫢M�d��3;M��j���4�xJiYw�����������������5�B��A�6�*!^P�g��Sv��{-��36QD	Di򶹖��[���-��R7ZJ$�k�c�0�nB_^�F��Jj�"�㥝��:0*�* ��n�̢� �P-�x�Gq�R(6�T��LV-R�Ef* .=O,i�;n��s<�f�٨�\��|W����2�K���Bo�y�.�u�Ȉ���T�����恂t�R4dj����-�9�5-��,
�R�
�$o8o3׼Ђ~�W�Vg��?�~H�|wpm�ݫj��b�Ov�)�3Q�y/gB]�QeMd�Ѭ�']]1��b
O�� �6C�U�;D������@A'\�[�<$�yGC�"T&�U/� �&���C�:�m�H�D�Z6�Ti�6�c�8Wݙ6hVE����(�;���i�����6�<aJ�F��w��*_���O��gCvM�5#�����%=�dH�xn�M�*ؐ�����"��Q?��m�0�m�l�HR0%���\)qm
U9�H��޵�|\�UڿO�`���+"��p����eig*�#�1�=o��b)!q�O�	���+�'�7��%����$H�����o~�զ]]�����̤��E���#<8���C;����ʭ�_��,*�#��Me� A�)J1��3����/�K};���,��p��*R&�/ڏ��(q���c�aw1���az��\��,B�����վ�Df8rj�V�A��:4�+Fa�AYt�d�:���ҟQ���L�����|�z������&�!ȷ%��|�I,E��WF�)���Q�r��$�H��7D�ћº$�k���_9÷M�����5Bj��1jY�'���ц��G�d>��AR�mnW�u�{{�-Cs؜,q�3�~��a��r��9l9��#�z���NO6X:W�p�U�ԍ��S��Hi���hV6�r���%@&���ll* �  ��:�2�ٔH	$�<���V�����O���f��K�0ykN�e��0=r k�,���Q�O�
E�K��)&�g� B�3��OO	sҖ�X~yH�t�ZW�N���a6	�Av�"����tg=�,��'.�蜗k>x��n�m��°�4�p�\��IR,�1�����?q�,͞`���:����ݺXz"�ci!DZ(�ϑ�޶;�"�y��K���B��P���1%EԦ�l�O��@c��X��?�2X�x�D�C\Tں��/�z� ��M/��nS�%�n��B<��|���1�ω�q�V
=�����{�l/l�-fǡT�f��5�{FO��)]���b��KΒ��[�4�X"�f:x5���X�J2�l��-hh�ʮiI�'x�O���M^&�>ǣ�S���Er�H��\�u�o����"R��St@?Ҝ<|�]�
���`[��JQV�6%t�+��=�I��ҽe�us�_8s�D�O,�ӓ)Ӭt��_��Q���"ĭ��uf :��Gnj�.�$R|�`�_L�*��2�P��(�fe��<��	��A�
U�&z��s�F8l��թ��HF�4|�^����W:�B+��S�_Yi���������e:��?��y&�o�`X!�ߍ|��6�M���� 㹨���d�)e_$��w{t�I~�K�=/m�;��W�mR�ff�����d�6�*�SE$��y%CYCF�nK^�E�������,��I�"����X[!���z����@ӵ�����<�m x���/�:2�r.i��6^ �����w@!���M/�D:�+w��^֯��1D��O$/���N�K��Vh�����z������bw���O�IE+���~�i�.���jZ&���%��a��#	��f|��O��CH��#�pBዄ���#���0imDF�lm�ՆnBy�iP9|���I�UT�/����\��ʅ�86�a,{9�2J�|��{tle�1Иס�2�#�x�]���X�J:!�c�*�0��_h�Ʈj+�x��W�hB�#d�M`�2 ؋��{/z�ߝ'�����⛰�! j����G�	7��-4y;E�y�2����|�E�`��b6T8�;ȫ�=�d���rHX��v��qy�p�J;�4�)����a��Y��*Ԍ� ݍM_���ٖ�L�@�w�h����`���N�TH�Q��������w
�kn�pAv���A}������Sءn�C����޼�{�2��vo�P�O3��Uh��U$�Ye�+3/A�I<OC�a�t����AORɚNF��.�%��W	�*�@ʿȼ!8���J;�v,��ӄ)qc*"�����Q�7l�H�a=�u9��Mb^&z0I�����Y���?�4���P��#��H���M�C�}�8�j��ެB��	�ReM|��k��xG/��_9��>���<R��8�n[.y޳1��n$�_����>m�v'�#�L��h��ut"#N?�,GX��
��g9�O�i���l�4u&�+��~��S�bl��V����86&d�H�(�I�D�S��U��\b���mQV^H%�t��́�ѡ%Fk^һ��i��{!�8�i������\$�'c������>@�1��`�UR��=�wxC	�4&j�Eٽꘕv�~��� i�H+e(-rK�=`�G���(�ˉ�k������TD"�Zw�S�Y��ȷf�7�.ج��Q���b������i�]��	��̓����Ss|��锠�����F	M�ݩUla�7h(WL�F߀bq�5�������|ExS�{��e^7*Y����-Ye�L���ݬ�8��9u���pcj�w�.A{��f�J5i[Z%ĩ�י/p嗍t3�Pe7�g&h�������t��밴V���O�'
np�V�S�
�����l�z"��3,
�P-���ЯHڎg�M}�W�2�܉2wN�ꝁgiO�O������ٜvP+:�=�!�P2@���	n��VN6�f�M���:���Xq%/V�$_C�W�P|�2M��8����x!�w*���:D:R�1꣤e9.=y[��P';l~w$�'��1K����{�&
؛����M�	�Y���P)P�}/��%s�J��uN8�$x��Xj�]�r�%�����\�����M��l��SM o}�3Eu�,��������|S-]"�+=�����z���CH*]9G~r}�Ę�M��Ӏ��&��h���$>��z����\�z~�b�M��;Cw�� f0�R9�	�]pNBe��U��Q����
��GWx�/��/��î�(�r����i�M��-<ޚ*�lA�4Q�O�:�ɞ��/�ǻ��v=���[��ş��>Ef���	�N>p3|B���>.>�R�7~[VmP���<m�b�sZ$�'�ֺ�N��̊����a���⇶��<�[8�j�g� ����d{�֡�+3�:�f�W�N
̲m�**�T	Pu��D���̑�:?�=fֳɑ���r��C�/�����s�M/�CD�À /��?j�����{�[mϷ�8�lop�=������l���S�QY�J��M1�>=�&�G�=��n��U�^5���K,��X�bEM�	U�����d�j-�EC��?�5B��.c�C��At嶷B�S�>��*�(C��ݝQ)$�n��X��?T<_�s�0�c{ ȳ�j���ʧ��tu��`�}ϱ��p_��({B�Y�a����T����i�a�k�C<�ʯԀ������{��)�R�{~�N �ER����^u«O�bMi����wK��4a�|�g���>
|�0Y?�A�L"o���)�wj�x��pd�|6�����D�T��;��
8da[(���]��_��<��V>��5�X׶>x@��	].��9i�t�:���s��<������i/X9OQT��B��=Wӟ�ܹd	� =�f?�Ml�Y�'1��%:23�r�)�N­����RA/����|�r������8�E�($�2faO��������3��#5���%V��pɵyeBrO�n�as~&���>��˴���۝�	���0��z˃o-��nAC��
!���/�cc���kҗ	�B�< OP�eA՜7ŧА�>o��8�Z
b$4�	2����0q�o�xDi�e9���T�vV���j��������`1J�j+�R�6���d��A����qԉƲ�3����9*X�ݐK��Y��M?0�vO�ll��Ǖ���d����B�p]�w�#j�u��p�4��j��8P�[�춞*G��`6�O�s+#C�J��4֖Mhi���)gp?�+��䅉�4�*D���]������S��
��
4��M��M�C��%�Pĳk>پ�&bjS�����^�OCr����]o�d����3�	Aˠz�5��,F�'��N�H
�S��k�<xd�^>G�>�*��"��
�g��!^�:w�0Q	L����؈ �(���L�o+��(��ԉ�����e:���z�%)����ȉڒ��v�"�I/�9����<����(���M��9y�%�) )U��p���f�1��jȁ��Zҏ�y��k����7�44�����E~��������0Μ�z�g'���+�h�w@g�uf�u7Fw�B�Z�]��hou>�QC]�\�eu��U�����1���u����>[L�6N�A+1��rq�;�Ӹ���$�׎O�}���-$�U�������xF���@��D��(it"��!�P����C��/����	v%΂��n�S�~���=�]Q;;�:�T;�3�C�D(�쳶a����-�E{:^-)�݁����	`��ٶ��T�^w��.½�'&pZ�B ��֝FsR0fS{�d��I�Lf������fB�UK�>��4��s�U˃0U"�&�-��b�V���v�~�L�(�C�岳q�ܱK�O�#�_�����/&;恒�YÐ�G��b�`�G��S���A��ԁ����|�r�|�����#L�c��I\!Ȕ�V�,�
��P���AjM��Y�Q�����e�˯��O�:�J�)A��U	�%ф���s0̳���j�O� Ε����Kdch5�|o�8���|�/)��W5-��^�\�AH�hJ�q��`�-�>�Iy1��sM�Q����nRޕ��j �l��;��ٱދ!���*y�6B�ڂ]��o)��ѡ�^�S�ͦ���m�t�k	vL`���H��+]�<�%�B,��%��H� �O"�N�L0�ed�H-�nr��\��?cJ"�������A�QSc-T��-��H38���	�p�=j>��¯ǟ��B\d���NŚXxV����,���7��YD�N�f�`bv��7!RAY�u���3 ���0�S�zd�d�H���ǌޮ�.;�n+��'Ix��Kf']�� ���n���dN���Q�%Em�$�w9�`�p��gO������~�����Gs��z2	Y�����}d+�rz�
Q���0�աTEN�.CŁO�/"N�)CfJ��L�v��WSf�!,db4MSp�}�U$����B�IxUUb�\&������ ���q�����n�{���gH�H�jN�l��A`GY��0��$��5�HE�Fq��;��zՂˍ���al0�vCv��^1h�7�+o?��]���
 ��\\��ej�4���K_��E�\0�M�}��S_&%	J;}�5_��gGOC��2��(����卽�/��3���,�|S}ٗBu�H�3?���G�C�FB<1^� �Y��Ԃ�"�����}�R�lѸ�R��t�C��ܐ��A`���f�p�%Ց�'�~���o��Z`�
�S���m��36�I�`(�79.�m ���qc�c���٬:rόբ� gU�՝U�Z-7cN��&$�X��=H��;Z;�i�E5�ƪz�	9�C�Z�w����p�(�wγqU����8�	Y]c����(�J��W?r
,�7O�U=@�����m��0�N�qj\�a���3mW�t/D�!]>��U$��#�v�:HX4B���(ӢE��Jo��+�\��>Ԯ�@��f�:[U:���/��$W��bEL�V���f������|6�$��l0>�;4��R��^�����9�k���<9�@f�f邀"�p�} ӓA"�y�34O}�����Q����j��.�pJ�b�l0�{�zǚ�vى���Aum;r �"�D��j�Dx<�'�>��r�܎m2��\���|��ʋ�Ywi�D`y.��$�q��F�W�[S�Ы���x�ѹ~�F�b���8yzR{�-��ԫ�{ �{�c�?��*��p|�� Q��Q��YwGZ�`mY@ Z[�@���e=^G/8!��<�%���0)��8��%�&2��W0\�OcB=  "�7eX�G=���.*h�O ���du����:�ӪJ��K��� ����攷}Y!g�[q��x���������~��u�dIn�(\�{�!�X5����]���a��ʷ�\�o��}J�0�]"��˳��H]���+ұ�qpo�/����r�pZz_���2�<T�^X��Mh�&릲@��>5T'=?0�Pi�Rm>s��+�F�s,]x��ƚe�)?�W���ZR�*J��T�0��|�:e�eă��ӚlM��DL�Ig���9�¼�)6"���C���{��C	rq�XC�%�gSC~'iG���g`���R����+�cia
�M`3�D�R��gj�m���zj�WU�����N���d-/$��p�Iz��ɝ-֗,fnx�P˔��%-�ۭ)C����v5�P+�<�X����#����4������&�C�KS�URtCUM�Ʒ�n!��s��C.��U�����D.�����Z�	�ip������Â��_^|����5�΅"vPH>�ú�?g~#k�-|�q>��һ�9Ì(��)���mQ��i��;�0���K������O�9�Z6H��_��pA���'�nn�<���@1�֔�Ľ����IP�Ĝ�������%p��;p ��L������N�dij�ʨx�Q��K�)�Z�
�p`QqT|[@���!�n�u��3B�ٺ��@1C�l��]��7Bի
�4����^�b?�~�D(��F�k���O�H�U۶�}O��*�	exiK�%IQLfLB��c� L=`�~<6�z�3� �3Kh���d�m���:�����BW a��c���K�eޓ�=���oU=>���}ܕ��ۀ�ށ�R����y�Xc�"t4:l[��{�Ӟ �
3��(��bA���5z24wv��8��:Kj�~=��罸��KY�����tm�3����Zv���ء��f�$O��B	~����䎨�z�^It�JJ-��B�!O�	�_�Y+�֮��q�֚�/�+ԋSo��`��s��rͳ�� N���By���jt}A�J4)��-6��C�x�ip�Pr�4jL6�佖�L�J�M~5��?_|%-�*N�d_�[,�|Z�NK����s�W�������o��ӂZ��fz[��m�\i�%�;ߕ!�鐯�ڡ��:rY����E�0�9ղ�Y�����@6���="��3����"6M��ܰ��2u��y��~3��V���g3/ً��Y�*��<���Uɸ�:0�fwt=��"���N��� �\)�
��m"T�#&T�Yt�3w��: ?*��
�mfB��i�,@��D��u�Sӆ��े�	�w������Z�mDL~��o +�uVU�6Yu��V�xm��fe�vú}Б�]K��+ƐZNY����Zk�^�r�� ��M��!n/�j��F��Rz�z{�&�u���q|t��B�VI��(�߅+_��+�2���"����j��J�]����oT����ҫN㖞4�!<}�����Ŭ���D-J�Q���am/fi�Ԅ����7�ڤv��~�W����9'ѵ��B�K��q����X���c(��^Osc�~W
�*&�g�7��g�)����"?����Y�S��̗Gf3��2:9:V�ZL�Z8��E�¦�F�#��awCѥ�+�M��6�a�^Gyis��(ѥ�4�	��h�6
;f��jț�PH5#��ܦ��I-�<�t<rw��E/%N�R<�D�"�2� ���u�{�p����gGb�Fgk_��\�U���ޔ�JǺW���'9�T�r��F�Y�r��C /���|���ѧ����,9�������s=+"����O�}��Z.��AwC%��w�?���[2=��T�+Ѡ�q n��-���Ht�|�%1����9ӹ���ǥ��y!�P�c�Mkje��}�����v&	�$�Z@�	2��
�m�����것�����Г�;���B8��ƺQ��Ɇ
�����u������<�O�;%���x�a �d7�F�R��S'���a0�k�{�b�t@	�"m���Y��/����.37�+�R	��(��� L� F��Ώ����dC���.c�Ą䶌�����H��	�vQ���4j R�¦ҲW�ޜlKXl���l|r9V+;�r��xK�ߖj��_��]$�t�7W
���/f���ʯ}��X�zi#z�*܂��8AT��+ZEGCTl�=ִ���r��[���ۋш g�����lJGƥ)Qe]��P�v����W��2�69�R��!�CL��� -"=���X���� �D��/���W�C"�eq29��e�5V2Î�7Ҵ�ƍ�}i'h�����$�w��4�tG��e�S�:��!��N�'o��:3N��7�$�fW0-�||���"�*�Bap��/fj<ZV��b� e�=-[,��1MVxK��Lu�W��[�$Hʄ�7JC�r�\��g�b���g]c��;�Ď�ɲ�D��B]��t*��x}^(@) ��V�������4�"&��M��- ԝ�1FIv�n�+ S�{��=�3&¦v�ၙi3yv�)��p�F�y�$��Υ��GC�F8�^*�]��杰��e�Anw� ��+��ɅJ\g'|�G�aJDYӭ����-��l�=7�"���A�~����[�ʍ�  !�N:�)=T��Lٮ�bb��ܠ�50�p�2���,����C7������➸A�-�w�'���%�ŁĖ�#W�^ڄU�t�ک���3~p�D���r�#ŝeK�lM��$��i]9R��CT0u.�����eK�+ʣ�O�KwA�S�y�*��������֋4�2i��ѿ1�����_�}ʸu���Jc���hV��ӵ���>��#�&��QJ��L���b@�҈E�S��40׀�Jr�g|���:/�ۋBTAɃh�nW��2�⭾��x-D�H���=�*:u+^�Q9S�s_�A�Sm��NGI[C�����h]��퉷��}O���?y�7T�7a�c�9�\�0�#TF���ZW�-��(�K�F9�Q�t�U���!�<���z �;���T���aPܱ�Xw>m@��ήt���F�����mZ.��6Y"C���� _锎��6R���Æ�Y��e�׽|�(Ц����=b�y�l���ǅ(�;�yqZ�<��D�Q*I٦�H�)������
;��bt�fwfT:R7�m:дy�����Wo��> 7r��:K*��n�Z��*_,�F�0e"�Pj��n�U�K4��*J����5�)��9*���������{eYU���I0�򳠶�SȐy�V_�������kaz2<��gC�r.��s��}S:�$C�b�p�����r8;�U��aQu~ @o^{N{�)dؚ?lk5j꟰+�qm�q�M��gկ����&�[nV[��k;��_S�8�zw����/F�����ӦCm�(0( �ֹp�{<;]�����������F�m�&a���S�Ҽ�#3��P��Y�W��ה�84�zu�0��H�w)�hE��{I�R�B��f��P9X��G79��9r=/��j��{�h=+a\e�q7@px����K0��˕;���%�,����W��K@>����0
(���N��P���l~���O�V� F���㌀sz۝��+-czc���Y�&S��9��a���m�c�)ƽGM��c�:P���4����U4�z9�+���ȖV_5m��d�^9Ꮻ�5�x���>�no`��")w�+A���f�m���Zx��Y�~��~�i����cpdJ�u���T�o�f�RS�ӭS�a1"y5<�["<<at���c��`�/W��HJ��nI�	M5�ˌO�� V�#��}���?��B�f �3A:�i��o^�����/��9�F�V��
�b�
7�I�ݦ34DΑ�fE��-b��q0�5�wj���x��%g���|���X}Ii�~�t���
�Ixޘo��&q�`�p����3J^JJ���я�-$��v�7�����gZcgD�V@ʣ�������Z�@G&�|��q^k�$�Q����܊�͂ذPp�L�ą���;��!���8�J�8z�H�tz��!�����ؑ.c�!���IP.U���6W����k��v�p���%�}�%Q�p�a$���=��ɔ�2w \C��숃=���~��F�����/��Bv�Hj1���|"���U'�S�)���k��$7�?���m|i�w#R	"���Ia"̽���Zz���B)���eC�ѐ�@��X��]-��N�p���0����0T玵\21�T��9��F'Ổ��:;�x51��_�xJM��������Uv���;��0�k��LH!<PA�RْD�-�8�|�J���o �5�i���"|���T@Z2�K��pNOR�s��)�XO��c6��l$��V�/�����|�n��@��oy��z厼��#�;�n��\/ '�E�+���uҏ��=G'ʦ�����l#Z~��.��*o�"Q��1����Q@�[>қ���s��R����=����q��!��e�<8�����F]����c0�_J�ȵ֚�`��� �5����KƪΘ��b���4)wLU�`�O��IS,��Ӳ�J���Q���L��`K��p�JWҡ���Tv�Ia�.�t�YB�NC�܊X�r��������v��P����MN�H���Mė����Ȣ(�����{�O� �UǢ8�7��F�%��YԮz0�-�|��B^M�2]�ƕ�>I~�2R��$�s��	/��-ݘE����4}�Q�}�Km��ۑb��d�:a�e�ض6�OE	��w�b0g#�Z)���m��$�U*�w�D�&��u7�wR������=[�9��w?����Ȁ
cXJ [����v1.9��%og!�rw%j�F��vۭ��BS�q�7ј=y1���2z�c#��EĈ�z�X����IC�#��ҋ�l臗�ݖ	���aT�F	b��|��l}@2p�zcA�4�'�s�<�?3�~pΡ�F�!��1�v����,�$g�˯a�����&��o����M�{���H�:�n&�C�*�\�u{[M�ۀ笈џ;�(�<���7�v����� ׊-����"^��p
���?��$��C���$;#����E�+#vl>[ ��:��W;��uq69�SL�/�o�H�ą�e�\tO�w�<��օ@<�g{n,�9 �`LH��K����PѸ)�#������$�s�`�ŨC�\8�����-2]�u��#/wv-���	7 &�>�
�ծh����G��th`�*���?����T��+g��W�q��f*z�}���UdVN��he�������K��/���ކ��k4���q��dwƊ���PUKO1풠qC�JJ��6x��}�N���>*Zc{�g4����p�|륐�	��q"g)�KӚ�x詞��,P��S����&��I����Ygመ oY�ܴ</�e����9#���2%9�.�M�o�`�pS]Μ'�:�I�!��	��~�=m��n��؟�K� ���7��a�ӝ��(c��&4JRe���(�K�D�GW���eJ�p��?3�A�e�ů� ���n��0)�C�е�g��Tw&vJ@�w����S��"&�iV�6�D/Ha-�Xhe�W������-��)Mp�T�,py�=���I	6-�������/�Ϯ�'�r��u�<z��m�NV�r���3Ð�ͤ��C�f�_�Ͼ�F�3q���t�A.�4eR�LP�I9�T�z���m��t�|(�Zc�5����/�4�-	�H�a��űz谑�J;�6jOS6�C�/��/�����`���"Y�s����4Úv95a^a���h�*�	C�*�\v�>V�7`I�Η���1�����tM��� n��Y-]��g���N�D�4�Px*�ۖn�I ve"D�a�d��B�B��	`H@�ũQjSq)�zĉ��U-��t*:[	�Ff��m�'k@������Y�����#n�?��#�I|��[���]�.���,ߐ�_i@��E�gI���k���]��.4�ˮ~��q��=/���cxo�)j�-�,�'[�����>�1-x�B�wP�8���u�n���D�|�6sFg�5dſ�P}'��@?�t�� !�0jV���g�l�Ƴ�F��7 <R/��ɘ��!�~[�u�޷��Sy� �9a>�1uRk�MI���YE,�9��>�'(b=YM3`7��N�I��5�'\�����R�E��矯]�p��c��Q�u'H����|����e�����qe�K�3x]�]aϑ��)e���~R����60���ٮ��٥��v6�����B�P��4H�Sx<
a�?#?H:�~��k�Z�
�����u<H��C	9#�
$xp�iW��jz���V��t�i�^m_��q*�<�VY-rk��~������	�zEq ����B��v�\��U_�u����͊�.0�J@�?�d�ޭ�ܷ��R�Wn=\�,�a��qO�u(��9N R�����r!��y�/�����<�?�Q����z�Cy��BM�!�X�m^�n��#����k��z]��pp:&���i/BN,w��^YJ��7݀�:D?~�,!=AK���ʥ�	��x�/�뗐MF�1M������]�M߲%�,��#~,���wX9��Oh5��p��,j���b�Xjn�>D=R_��M�TKX4�}Z��	��"k�|x�
>��j��h�T��N( 'p�~�Ps�ZY͚���� 004���_̄�<(�ܔ� ���p���������a3��V�Gg.B�&�ȊO&}p$��z��~i{�JX�p��}��ϟE��/=�;���iɌ)2Vn�.�TD�D/�0�8H�5�[ޚ���Jwn؅1��7QN_p=��ߢ�#��5�c)�0ٿ�ˠ�\t��?�%�6���r� uMع��K��F[<����������^��x���pgf9r�o������I�_��}�Ժ���D�����J��R�΀$AC>�"���\֊!����Q������l]MLC�?'�K?4��?�=�	5ke��\�"�j�Hs�ب��;��_��QR4���C&��;�	f�,�6Vm� �P峨��b:'�%3��>�vR�Dejټ����gjM��~��*9���L>�WF�q�׶�Cg�K���_���a�W
��I̜�9~�?W"o�W�)��1Ŵ[�N<iң�6���6��#����w&�A}.~M������,s�qD�K �\0�%]� ��E���j��~8"8��#H�|�(�W�S�P��T���-��M�KH��[�T����lRd�WP�	, )����}V��s�w��C��5���δ�@�m���a�@��)� e�%c��$�[�����)�n�M����S��gDymx�	7q<'!g��4¥+k��J�s�LM�نCʄw8�8#3p	�E^�і�T��� 򅍻�o���#�-<���:[�'m��:�r�tdG�������kHd�j  ��o��`�?�+s���B$e9`5�p���
���F'7�w�� {���|V�a�"1r�|Ɵc�m���`:�௲�]@ni�`�a9:��[��.o
��lٰXg{}NT��X���m�p��z��6�GQ�!�N���
u<+��XW�����?���]����Y�iE猌�Ս��[�*�-��"�@,U���P��Hll�:WN��E���.l���?i[^ꚵ~:���t�MJ^n���6�I	Ei؏�V;h/��Q�z��2�,��U��rJ�˵��{s-
�,kX���9�J��m]�Ը%�,�>IA��T�5�d�$�3�������_9 ��p�;ՒYQA U_ʿ3`��1�9o�`��T��
����ef	�y��[�G�=�Q�L��{�?�K��N���xos��j�������l&x���W��*�vT&Dq�,}��i�婬Q>U�<W�ƩmZF�(\<r�o���R���E���K�����CX=wkr7�h3�o���U�n-Gr�=�U�f��I�m��h�G&��Mɕ�ƅ���ɥ>�L/�������}�8�����;*�/k�~R���ˍ�"f�=����8`��UZ������>ll$��R�n;L��b�nv�	���o��dB^RפL�!��!�G��$ei��J���M�)^<�t�S*4.4�j����R�s���4�>����@���g4�j-����Fjڣ�>Au0�@;����	�	`ո��B��'0n�ӄ�#9��R۹iQ�(�^��46���F�T2Ga�͘/��8�y�	S_."���Q�DZ��h��`�A�����@x/��5?�X
:��q6�<�	���ƛD��E��FcٝX*�&Sj�X�í_x/��4|9�pu]x<�)��W�L�sg~��8�K/Pʁ���Vf=�6�#��3|�&�1/gd@�m��pDP��y40KD%ۣD���V���������rFɶRX��b�]N���P
�2a���-	�`Ζˡ��� Me�[�{/�+Y����kv�3(�B5�'�d�"��O���i��tci}�ӚF�/X�褌��*�	��e֭p�I+)�,>��+��vW��G�J+�1{N=�r��_��!+���ܞ�¼�*���N ����ia+>@���s���]�s������b����O���L�6b��0�d~z�GbG;�ٲ�%��������gVO��r��&Hp���ð� ���X`!�鴛N7�A��ne�����J��ݐ�qfnP��s . 9�a��G�Y��ulJ�	��6��dw�H�w]Bک�~�Ȏj%��.�+��ݽ���:,�$ڨ8�\e�6�-�H@��2�{&~��q:Ɖ�5�w������7�o)�_R|b�&k+j0�z�a(�M%7ѿP��ETv-�j�xߗ�$�m��������"	�e/ßXGU�.?z�W�N.,ߔ!��6�Ⱥmc ����S�/M U���M�L;����e ͇	��M�[0cN��&�5lFתjW%ɼ1��f����j� �Pp���`;�C�w��*��V$9��_��� �.& �q��XB�TuPY�cV��|����8�-��ˬ�����s���	��6�6A��2�%3���<�]�{��`�&��g��_]�`#��5�J����$��Y~����?͂uw R�|.�iH��p�>�Ih�9�ԙ�+�����l�շ��ᝪ�Z���'@��-2]*ǐ��d��ΰ̲mׄ���g8 �����m9�$1����q3�����c�Uu.����HܘƯ*7{��a=����*ؗ�.W}�T��k[j���WC�n���@x�eiH�^�98�==�~����0�u�Ƕa�C]�-��P������},#K�D,j;��=j�=$����tvY]?�������Uc����Z�#����M��^ŗ�2o�|�71@#=2�ӫ�<���~���+� U���,��R]���J�͠n�mw{m�D��S�7�q'!��p���{��cC�����Q��1 �}-�7��ɦ(�V_�?]�X-�q����&����a�R��U��P{�֛�l�^�qjlH�s�������ktD��g�������,�c�M�g]�x#�f9��S����Rz��V%��A��u\�V�֦�N<�Xb�[���LJ���_W�k����Ql���������-���X��W�4/����5��T�~�Sx�&K����3�}d=�;�OA�OB�i����=�b�Hՙ�sbHtkHU�'�{��<�x�\�{��R��Crp�rE�kp�s�{��xs��DO��aBƩVz�5if���h�>�8��j/�#�;t[`�r�1���,	Z�Ű`��ȴ�'j�OI8�?��e���gU�q������f�貇$��N���a��dg��w�-���MflXx;9^����Kv��V���@,�c���'8{�z�����%�@��C��x�%���fێ��m�Ý�w\�RL��Ȃ��G.��6���*G�U]'2y�5����g��X�|�/L�\8��jT�ڏ�-zZeɋ���|H�ᅗ>����#Y�<$�镥�������xA��al�P��q��U���8�B�m��B!�̡�ڂC#�׳n+�|�HA	Ma��ig����]|�ۉ��E
]���_T�M{D�ƴ?�X�ԭ����r����\���sK�'�Q\�և�X�l,�[$oII-䝒�@.��o""\�o�?�,|��I+�ƨ�S���:�6@�a�IG��J���H@3&vb-�緭w��L���,w�*�?zk7�z����>�?�φ�����
��-�J�N�9Z����zsl4W���zp\�����7Z�d�Q�0�.]�kZJz�����̪*{uI�o�Ɂql#�;��&uZ/�ZX�\��<GTc#�k�E�/�י��5fS���mFV�A�8%d���D���*�����־B�;|�Ͳuh"TK�P8nt��Qu��k����a��yE�L���lŭ���;Q�4��KNK�|�{.⦫�F~q�u�pm%������ʹH�%������,'S��ÉK`t�̼��yp�\�z��ׯJ�DS��WZ�Y�ˑ	�3�vȷ �@�q��q��<�x��0T�S���AjS�NC�����Nz�/�L��b���9�Gd3�h^B�"��5S*_n���w���s����#k�YN+����>�?��e 3q)�4Sӗ������F���b�vY<3��2� �"�_�Ŗ��������p)��Wl;h�\� V��G�1��s���ĳR�:��ʾyjl����^�;�Qn�� ���XB���p�`�4�Yj'G����::�Q*�vT�<A6C E�Ȍ�����r@���$���y�P����/:
ë@}���Y�#il��--�Ky�U�f�6L�;5��j>Pi(���zr�(����������P)|U@�d�;$s�Y�dE����ʀm�|j�:��=�^!�|j��t�����c�T�B_�
�U�?�elЭ*6�;���v0�$�#%���������7��J��f8����_���ɟ����m���-@z��<� �R�[.�H8�P��]@��m�ô�g�a?2r1���9Q�Q�����p��A6��ܦ���Zh�c�ٖ҄��d�`�tmK�&�Ų���q�){����{�h��̧	콒i��;E�;鉍X�uz�L��
'Ӧ,�<�\Ň��j�<��t�o�'Sp{�>�Yxv��E����"d��(�OYm��\y>�^N�� )&������SNL⠇^ޑFd%@L��k�^$���k��^}�WPh��X�F��뚉�r� 4���'/���ڸ'�Og���гNVBl0��ܱ���Nܭ
)j�r�MGY�Z�;��Y��������f&1&$���hSSqX���k���_�U�3p�;p����
f�%Jj���]��2���B��z���9݊��̐B춭Tv�I��xR�|�/9��R�R�m��S]�ս/��Kbj����zF���z>������md��޽ �?3�bC�onIݱ+?X=��3V�����'i�^d�1����gsa�(*����U��w[�x6��[�\�9�
�v�N�U&����g	M��Y1~�kBt��#��zƀΐ)�����P���IBFM5�m_�i��h�8)�I߬rYs�A"�ߺ�����A6��* ����h�{��$�$�i���w[�i�DA;��XF������_¤���� t�W/øF@\����E*)9������R��
%�	$�R�|%��,[��*OB��À����U�yj�W�`x}�6�I�l����U�p��	�!���	��e��z�){���c����*�ٲG�Cl."Ѫ|�T�@'zE5_���)��(��?�f<���{�K����IF%Z���k��~�&�`��~84d��M��*dj�K���t�['� 8m�h�*�F:�M����Pd�]'QGՓ� �0���=(��+���](�L0��[y�#Tw�g=�W�Е}*)��}N7�}�Fm��V��c�e&�-�m�R�|S��VrQ�l�a4b�=�����4J�X�*0�&Z�5]����;Ե�<�^�I��������ǐ�߻K$������~�h��C�OK �l�ҙ�g�������6@W���k�r��YFE����ɛ��W�4�y`��G�n� T+���v�j�UT:$���>�MDn�^���덭�B�Y���@��i'�:B[�v�`U|��z���Q�g�IM�O�?0W�v�P1y��`�(�f�>�Z�qJs�3�l���$è\Q5˙O%+<��[W���2�N��Ww���&׭�b3G�*Γ�A��&"�jv��П�/�G)�����R+�Q�M�`�T�}f�`5dB]C0i%Fܦ@��ʬ\HC���Q�0�����5oMh�h�n��k鸌����{�)�!K���ДK�YN�zC�j���@�я37��?T��K3\���-:f�9df���7�AD�Gߣ�#��,����#�@aK8�1����;Qr��ʜ5�����Pu��5�CȥN1��Y�[6t��L5'e�U2^��զ���R��4�/�g"�CP����S�@a��}WDD�[�ta<8�D��%��%��Iv�6P1���h���W�B�q�w,�[	��'��@�P�w����D��-QW"�gg�$}x�DB�U�����ōx|d�P�Jr�Q����q}�q���O�ʍu!Z�,�����(����:r Hx�!�hy�L"��Z*��rMkd�������p�H��9�q�t��¹ŠSL7� Qv�j�_1�B~$�2�(w��^�n��Y����l����h�Qek�<!�b$�t���'���1�H�D`���x�%n�Ü5>�ͥ�dϵMb�[�1�K�<� 4��@��Xk�A���-~�L� ��+ m�����-E���GQu��2��zF8����d��09�p�>�W ��rj��{H��~m�|�'����+윤�MdU���T���hƉ\�[75W��♾/�=�&N�t�n�{鯐�qn���I�F�h�Y�{��u\HzX8��ܙ�����>Fd�M&wh�½]�o���@��F�w��S�L�%MYg�f����,�v ���D�4��ɷezu�0�������	^7#��z�,�J�����(��4>zIJ;��)�4ط4�+��lm���S�r�a=	pH]�GRF��h���[U�h�k��`��{0Z��Rݔ�&H�/��槽�}PL5����ջ�۷F$�\�vT�Lm����1��+O�c��s�T�Ɂ����'&2MKʹv�ף;��~=+��#A'�練�B�d�8~��Y�rǀW�*�*NnM��qX�&����?��]ZbS8��¥�=�1"(�]�����krюm�3�5	ma�0�8<�N	��YD�X��xLf��=��л`��)�+�RN���
q�?,�%Tb�Э�XBk�=T��c|ok)aZ_l�~L���<�7�³9B;�n���ë��hOS4b{�5|TV�a�Vi��h�zO���x}WG�R���z%|�̝�y����a|H�^��/��<3�� �֫�������0]JtH�|a�f��ϟh�J�`1�6�d�4b��1��!��8=1P����>���Pzk����Hs�"Ox��S�u�J��d2�|'�����PR���C-e7������X�n�C>����b��ۭ�Y<�a3q��~�`'~W�
�0]P�B2��`	ˆ���\�p��T���׆�s��R�Ӑ�_R�X��5��7J�:��7x֍2bS}Q�W�V �X�"��_b�����V����E�g��Ѻ�Y'8�3����5��y��ZB?*ށ�晼�0p)��L�ưur������jq��)�H� $[�m��]�~��0h�^�� fv�>�����y�~�;N"��-��!��U6��c�����/�Y��0�k�eͭ)�N���ϵ����]�7�m�X�_���w@�("�%�e!�q56����q�_�9�
�2&��
b_W��C_�VtQ�#=���z\(QN��.3�v�Tϔ�W�&�����dDH�FU�{B�K_����4�*����÷��-mw�fX��.6�X����6�`����7~��Ix7�۫��%�7�1NRg�1N2B�`�&sߥ�t[q���5*�\P�x��Ŝ�̟K 6D_C�3>بJ��ww��V��|?���/��B�a@�t���f�̓?�Hа��ec��R��9�>��׀�%����(;JC{fpc���g�d��OG���0 VYi��2�v#��Lx�x�d�e�O���0e~�	���zZnm<��D��*��pG<N$��z7]ܕT&&�^e�x�۳��b�W��IV�&\��#}�����?�u�y�J����-&s.p�4)����i1���l��5B�4�����>j�\�\���=E�
���c9����#�7�y:��co
�>y��J�.)!�Y u�%q���������[r����(�&�,Sc�8�4�"���|fU�pB���v�=f�N�0���-�Ҫ��gǃY`
9�
�d�6�HS�MV���`�����(�i�ow�bP��������`�"WhL2V{b�^|�>�u�/<F-N��e�v��d�-����f�Z�Y�kU�힦��k_�b��ѳC�����l2�%�vr��愞r��!91��E�"��9Q�6�vZ�'Z�N��P]�e.�M�j,KE�s�N�W6x�3.)0��_�L ��v^�9œ05;S�D��z�q�V�7��]�Dy�.����r���Bd$_S]�����e�N��<Uj��\�� ԺRN[��?yu{�`�;V`�T���5wD5��°�g�73�`�u��ٸ'St��I��:j�4G`����s�G0̝g=���}/N���,?�Ń��bWLM"h��y���w�vp��/���W��C���\�ht�(�� ��oY�?S�3���1�?���V[����,����?0	��}%�}9�	{e��
ZS(N�=T�Яp'�?Z(�l�N���߀�	cs(n0����_���д������7ǅ���pVH�ZdyZb��<�z_N��X׿si40ZW�bO^<���6�g���N��M�>N[�G�W�h��.�T(A;�(��#�(8o�	2�`մQM�Q��ޣ'��X/��딂�~��~꘹zc��b7
U2�E�@4�mW��u�-�� ~9B=��^D�x
p��#�F�B�y6�7-�W$�S_�.���y'M�h1?����Q����!�ܘ+��
]4mmZ��6A�z�;���ix�K�:g�в
b��R���Ȗ���8��YE?�M�4rK$/�LU�Ά�KW|(�Q*�4NZ��<ext4��n2���n�*��D�u��v
�u5(LN�X��aRn�(�pF0'�~UB�1G�0�3
��OY$M4!?���
7{M����Y+��r����"�8���P�1�־V�_;10�VI#�j��F�@h:����!�_�YO�*tO�C���{�4X���oH�4o�w�E���ѹԳ�5�Մg��^��.��(Xk�('��I~���D̈^
���rp��8���%�<����E�h���#F�L�q̇��V���AX�)mSb��C� )�4��O�3�S��_��})���$�=c-��Bs��r�Q���`�K��rK�/�@Y���������Ч���N>�N>��僲P�-[Sw�f��kuN8\�X�r ���PN���f��&Z��� ���I�7:���^'*����	�5���LSݐw��~n 8�WroNHk��8�\�8(�M��T�$���=_f��� i2l�Xb���;Ur��Lv�Ҹ� ����;RV��~ʈ$��?6h �P�|Ӯ�e�b�Z��H�Qȸڎx�?ntiDSMH���S_���!�z@�,4ގ�/��تed�-e|�����1s���q�<:/�=�}��Y��S��rL�Lr���X��,�7"���RER�˷R��|d����fP�@�I��I=�r�3O����%�q�KQ���%{��<.�g6@7
yu7s�h�j�wZ��0�i�ɤL���.a�9x�2hv@�'L���%�ơc����s#�/���U3���;g�~�;��ꬕ�9��(H>:�6�sw�U��jGB���C5ޕ�U�.ΩF~9D%�e�@4�ф7Ī�U��0��S�\��lR9T����N�W_�܃�T�֊�3�T��V���b��OzQ��T8�?f�ne��Z����U�� ��q�oY4�`:��8�^Zv�?�����p��#{	�e����/��h���p��nH	��M���|,�Q�G�;�?/Q�:��7���i��A�X��H%�����;�Q�] m.H�'�s�k���q�\k\X��uǔ�}o`�K�+Ks�yyw_���x@��1���Ӟ>	��'��N3��7��,�$���3�:�(Dr��sQ՜k�K��,��n�	��œI�M�ً��$�Y�5.��Wa�h(9r6�g������PM���/��Ʋ��y���8�&�O~T��UJ�_$�}�qz�)�0�<F	}{j�>���_�0�~8%í��|��Z���k�?�)\J�����&˾H1��Bo�b��]��C*�?��������Ө��v�X��5* �1Kv0z��{--E�H�:+b	�6�5�E2�����/�#���e���֊�vbW~����_�&.k��=~�*ߤ�1���AJ��Mώ|s��k�b*���|V�t�?��Nݣ��y���h����*��߭���N�9�����kԼ8*��"`r��Td�g��8u}[Z7ӻNW(~�~�؏�̽}����[���A
wDRT]��,&��E~L)�r
��<C�pc��I� "v�m���>�uV"��q���ijBd��-�q�u��+����̖Ji�xar��N�a[��17�/��`����2Z��L��?6�p�����ힸK��J��nȗ�^��}#&[�~,�a^E4�9�P��z؎hn4���-F�8ʏ�6�v�Bmj�?'t��yq�_~���^�� O����l`�Qnk��r�����O�ܱ+����-_ḣI�J;M��-�i*w`?���=�������\��)1�۾�Q~�?Z��|M���R|Y��Qԉ(���J<��>��=�+aS)C#�m�O4��RJ�S�r�f�I�(|>ei���ݲ������z՚�Ħ��g������dc�o�MȘ�S'�U���9du�����n��^�J{G��uH��X�#�J7�o~�R~�(m�m0j|��='QT��T����n��C=U�-΄[��!V��HҚ�hu� K�t͢���%%������ �%깹r%�L�~o��F
aH����H��������^��B(|J��#|��7׻��y�5���	�� X��������g*��e>�C@��M���/���(܆��h���Cg��`i8�O�[��M��)"O�!ǅ/���tH�(}]B՜|�j��S|+ǋc&fX��1�~��n/jg�8z��
�t4Qm�υ���()�����aߦ��ե�῝����u�$Q����M������~���+��z�N��~��wh�m�2ǐA�/<á9R�.9T橪:�;�E�RU�szQ�CU�H^\��Ext�V�5ʊ�>Ym�6����f��:3;Ķ�i�^�YC6׃�O�(�Z�����{磲!L\Z4g��U3�nf���s��b~�&�T��TNTr1=�m	ݳ������K�<?�j�m�������hhe���q2����D>��%�h�	�u��J赳a�������')(�-4�y%���/�K�=���b}�٢��ַ��V��<bP�kԴ �?W��S#�17+Ч��D���;��Ձ�/ચ���[�E��:�3�t����H
�v��8�QRweq�<���Q����
J��q���?n?�0���X�$z�4ɝ���n��:c�2"��91<�ό�rZ6��y?&�f�)7w{(Sĝ;�m��)R��8���FY���{~�3�u8�w��ÿ�w���3���2,���V�r��-	���`��|�L��эtQ���ߩ#G�>�.6���h�Ӟ��?"�ol���/�jI��OՂ����Ooi��aV���T�!,w=��j��K�.��.6����磥M���O��H�؋�_���r1YB�J�!j�����i�8i��?�
5-�i�%�)�W�X4��]�Z� �2��)o��w[j��cwG���`?���z:~�� �T�~۟�O��@�o�߫�I]�~�{�/;��P����m�	��{D�����$5OB��m��N���11����O�wjB�~�U|;�0�3��
��ceL$т^�ϑ5&sFM��k�'b��\U;��!H3bg� �Zk�FL�$�d"Eז�+���Gn�,�b��#�d5/�U]t���.|$̞ܚ	K��X0l=�q�&A(B�EL?B~Nd�t������^�L^�x~���4t��捀�ϐ{I��V��E�q�Wb��b�[����@!�� 5nZ�S�1�̇�W����-��
���P�9/fm,�Bd��Çwj_yI�cue\nvjN(<���v8����l���,R��2q����~�v���ǃ������ƨV������,~����e�����X'�:t�]HPYT����ҥ& 7�`�LW��/��J�T��n�>����̻���Fy���8��쩬��p��v2�8E���|P=�	�f�0PIV3��OQ^�*Ǔ'T�>1S�Z�l�~<q�X�΋b=�%]����/���<�.�wJa.*��{�ӊ�S�:��ִ��6����FB'o�]N����u�'�,��K~�E���{�N��4c����S�fg�JHe�U(TKmԅ �q�O�z@p��#��7Miܽ�����nh=��A�����p ��TE�5�?�'��G
�_P�� ��f�-B..	g�#�x�{���!䢴AL�ct��lV�J�&>XSYkeb�f8�=M��5�Lr���G�}��1-�~��[�o�0B������]ϳ�����>��lp����o������ sV�$l�T�_�!�х�fΣD2��z�9�� D�#��^S���E��m����vY����+-��]���2k�0�q����V����_H�_��8�:g��T��nH�{����-�����Mt�-yG��iH�[�L������$4���F�&Fx��:�lC�d�ڻ�i�j�J�����{;[(���������f��U�N!�^?�F�%�nR/�?C�v[.��F����<��M��=#�CG;�V����9��Ǉ��K'c��5��̹��5����A_�t�,��ґ���r:���.{}��R��E8\��\ŦE��x#]�k�AE2�(��>0���lZ"蕏o[�Y�6ni6r��� ��vc|	mG�>�r���^���u��NH�of�d�������':?O���5`�����o3�ϝ�A 7��a��v�.X0�L����♉�o$[���Ϲ�i8I�ۃ����&��K���q$��	j����0�2O�y�a˹8�h�^��I�#�h�����MWH�NV��ys����2�R�c�V\���9x�C�2�[�/Z猺���#��>t�ts%R����u�ev��q�e�U�M�o[ajȐ2�3�5�4�/��>m�JXh��_ݲ4��F(W���n���4�,������,�"&�q�x@��D1��^.�u[
�vbd�	�ZׅڧhbFN��yv�	8���Lk�4,/8���Y�5�Y.:is�����]��!�u�:dB"T��!�(�e ��
�=Y�d�Hs�^I &��~_r��B�A�.R|s���ښG'��8���o��A��2PG��^
����t�%]s�]8j�UD��C���p�O"�7mUy�������V�D�����6�H�cu���=L��n�ܬ�!��g�e@���z1=ܠd���^̜[ G;�oĴ�J5��s)J�xb��2���h�$ft�:
��y�t����z`�3Y]�d�i������>��jR|x@Nd����1�����R�=B��K�Zв��5j[�Ɩǉ��5����g�SJݴ�%X�:�j��	��?WS/�-N9z�G������;�p84NcZſ^�{�B��VĩT�����G�\7ɴϺqV�U������W�Q~��n&��Y�HC���ZvbW24KL{�	�L�05�b�v�q2!lt���	�Uk
~oXW�0��R{�|i~� ��#9a*�;i�V t�)�oh
�u�	4�������N�^[R�z�k8C$�
�:�V�F���Ş��mx	��o���̤�hE=�d�$(:E���a�uo�$�m&O:�� �`�����Zw���6s�|���i��~gȯ9���u�Զ��14Ӈa�x]��;�m�����AJbS/j9˜@b���1f��0��j:
��$b�#q�ݬ)"ٖ���Ne��=C"��o��U, LA��&�׍��cN�v+������T���:�Y�ۊ�d��u�5�{l�$h9"��@�
U �Y9��"�'n�l7�d!�5�&�$��x[�BF�KU��m�#�?��}�#wo+�f����J���R,7L����N���_�G`��S�&E�C������}��;�E3E%��ŋ|a������
&*<PEi�E��#t��C�Mt���N��*D3z�GH��G�{��U�mD�-�$D/Ò�?�$�"��i�7<g�N��@��;[�ׅ�Э,D"���Y�7��R�|c;,�T�'Kij��c{�͐�k˕W*��ܯ�ky�C�	L�!�^��)������?줎�?-���]���I
i�%��89,p��D���vS��o��X��NV��cO��k���+�)/�2�(u�s����a��e��"r�U6:~Q�0��
�m��3�����+�Ȼ����y ���p���V�`'_;mh�<��ż�>b��r�ԧ�"�-�-B^^���������&u�B%��r<���U�n�Q�Xd���P�ܼF#���TSP9$�3@Pp�\*�'����=����35� �Y&�L���ܰ�� ��y����LX���!�џ�����fz��0�Fһ�ǫ� ���Ox�6�b���=hQ(͆9/�t%j��(%������n�n�5Lx}��� �A���3Fɽ�U�npWl��@��>ɡdR���b����,�;��C���8���|�-C?�N^��c��r��5���e+���M��)�p��F���lOJ����p�L�h�;_��)�{D�m���d��7/S|/Vf��|��vIJ8}��:�裂�9���~��oȝ@BLz<N��F'\�/����Ƞ9��s=�9��"�M`���G����3髖��L	��ѯ�=a���Q��Q�{��7�v�+��k_���M�;
ܭ���[��C�0t���Ԩ�A!�Q*��e{�07<~��-���+QF���+_U9�8�������<��Tj�nS�����E���E�%,�_��k�|)�p���SF����ْ"X��?����[���Y���MH���ev�YÚ ���wFqY������+��+�,�i�jC�8�8�Ti��D��	�[�\�d���ROa�42�6��C(t*|���P�����ߋ2m&�j�s�T�(S�Ƕ��4��0��b�U��L_u ����~[�x�zI7��dڦxV���� F�~L��h 6t���6��t��Ӆ;����ŊO���S��#�)��$4z�l�50�\	�0&����\�d�����u��ZO|�@�� z�Ҫ⯔%M��;�^9�E��_,�@ӨA��B�9�� @�/�'�����|���r���ԟ�ۘ�XF�{����v�B�$���$g��C<މ�/�o����,4��\���hu���~�|^�hk����q�{���?�����n��	@�Sj�˯���$|Dc���tb���w�s̐P4@��	�xn�{�����I�C=�/W�\�����E��bM��Y'�JF^�K����L�� o�BS�t���Z��P�=�MQ��t�p1��7��� �2���.�8�ֱL �E�=���R��n\�3���ȏH�i� u�]Y�R�w߱y��Fn�p�����rk!�w���R�g���|��^�O��;������M�*0��Me2�b�,|zA�s&�y�0j�"�#��+zÿ�1=����x�^z:0$���TG��]��[Dp��r��0�� �d�0�(/S�L�4�'�A/�r�lR��v��&k�P��a���g�>�o��3 �k0m[�H{���s6`�*~U➒F������c��u�a��c�p)�THg��6��CV�u���_-`��d)��Xxs����1�w���OT!RT��������k~���V����/t?k.�;�Ũ��'��81[���3r$�_�K(�D[o�]'I4�E�+X����Q��]�2�T%4�� P-���!fQ�0p��`�O���n-ڥ�����i9> �&�:��6��#�Ohom-��)�'V$�/�3{�	.���-9fՂ�h-l>"��i �"�X��9]_r��䶴��	���ç�M>l/�%���n.g���c��4w��.]A��VF�e�[g���+��>|�I��|�������ԥ����w/{+���	��|��B����iu����`�ÃER �H�(����eۮ�4R����c�B��UW �:w����F�M>Q4��>�h����	�+qk�piDW�U!�vƿ�z!�ɇ���RB�w�5�z��!rk���Z���ن��uz�j_j��ք=ç;r�r�q"T�����<"�М��H�}6ڊ_�e�'7�tE|F�WX������"���ɠx��T�.!"�c~�8��k��o�����Ii����� ��{��$ݝP��L�d�R�}�� &�{Ƃ����%�r^�wc��
[J��5�Ș�a}'�+�;���ͭ��+�ň<����mgs��d�;UG���'˭�W�Rb�4Sj ��1�Rۆ�q�P�b��_�I�u�����]���z�n��Ռ��K*\�V��m�� �|ԉ���&ްY[��\����ձ������A�ʠ��זy���v�u^��!a�"��c/) '�	A� >�����!9�����Oծ�d�E���)�^�*~E)��-��݉���o8�{ S���3g���`�'�L��"��wvc�8d��v>)��Є����W�H =v�^�	HĬ�� ���[|j4�Kz	�%2����"�띻��PX� ��S�A�j쀙�`����pvb/��V\b@n��ݓ�k`�����	%�෮�}��I�	XbBaf���G�Tͮ4�V)��֕lD��)5�R�F��J�
μː�
]:��@goW\|�F��0�K��#2c!�?Tm�wd앩�;�*?�
>~�䖷�e��O�����i�GG"���f��;KS�U��$�{����K�� �J��Q�J���iy*(�*7��9�����	$������K'r̜�-n��C�G,���L��K����[ȸ�_�X�k쉙MF14����
�鈅��"�p�d����_U!���Y��cm�؀~�k�jԤ0��9��N�ߚL�&,:���˨�v,���b��;��]�����^#ծ�b"�n5�/��L�g��m8Mwt(���A_x�
L��������F�q���a%�d�c��("�3ͩcϘۂ}�d���)�n��ulGM��	XD��+4�K���]��՚Z�� ��ä�;���2s�^��+V��6W��O:/����'�T���[`q��5Q�B1"��}���(��N-���A�v��ȉ�-�G��ؘ׼�o8�t`2s����v2A��R�\�\$��g /�޲�6]C�ΐO���(3�~$*�s������@fZ7f���6���N"I#��J�_��0�b�_���-���}��"�(�N�e���>x����)�.����삥�����4X��a���~���7����\���+$�mq��˛y{���#-u!��9�Qn���g�YXhkn�i�<S��������U�U�P�7�g|�K=�6�GkB��V"��n����jz�6��ҏ�I�Vy�`�0:���8�I�;ZܪWTqV^��q�����-�ה8�#��o��a���g�� 4��ӆ�*�,S�"͢����_��,�6��tj�n�z�ϓB�XY'b����0Zu{B5�D�fE!�IM9��|�$�_X��UA��td�ޜ����f̍B�j@��d9{o���[,а���#���ё�"�@5���@Y�M����=�%�e���I��d��ly�3B��j�."��4t�Y߷�x_�ȴu* ����c	�V,~�_8�ż=��nx��E���d�\:Oj�G�_f�;@}��a�Rq��F�����.��{r$b<�T��-��ueŒ�+�:2�95'p�#��	~��S6x�]���t��dv��N�|˸B��-�����w��ij�i�?��<�h*�j��ߩK�$i�S�6�Q��t�U_œ�!.马gHґYmOf�8ý���U��I���tXM>��9��'�Ct瘲��Md�܌��q7���9��[ʝv��UM$�e��-�&ԃA.FO�t�Y���: �/��E�(e�s������4��!�'���kj��/�+3C5�S�U���v�^l����MR��PM/���a�ρg�|:��"��y��3ͷt�Q_��F�6"25j�$�ad�k�L �gkP�Gl�ወ���T�M�\�X�	|��$gN��HP���_H�B��R�K<�-u!��O"�	ìw�A�KM�4kЯM,�F�-��&Нk%��
�� ƫ�����M�����&J�I�ކeO���Ƌ�mm�m�������E ����� =�`|�'om���~H&sB�Iu%!��P���6?ж�h1Y\��%)�D�`���N!ޘ���\�i��}5�5T�rpX����m�=������e�P��>�3�aῳ-᧫�4�cz��F���<�v�����>c�*D�{�{f'豹��pIx�EgN�T7�_�����2j��A>W[�xi��Yx�P##!/�*Q���d���G���H�������i�t֋7f�0TvבM���Ⱦp�jvECĀ��p��8Cјm;�@i��Wpa�����{/ynz�gC���Ջ��Y�@aHM��ȸ�g��tUJ4b��8���$iݖ�=��J$�|\~.�Y-��4�Ӻ�1|�,�\v�݄OV�p�ܓ|q���ytV}}�ތP]��$@�zzeZ���R|���b�d5������|j#ԟdc$����aL������^^��e0|a00���|0�v�`-��A���A����E(,N!�0��g�����4��xO�w��z�dj�N���a��W�2��_�� �=�I�#�i5)��I�>M���NX��&>8�..�$"��`��)��%��̘����Q�2C/�뵻���+.5f�O/�e1�i�6�[�c�s���Z�U�\�F�o����V.Pk����.�Y�,z�?��y؅����i�;����h���|���k7P4oB~�Wi�{�?�R��Fn�aq���?#aƉv�PY(L�~�a#b��]#�:�y�rP>�~v*x5��Q����!mS�<K��c(UO�ؓ)wXOo���I��j  :HON��g*X� @@Py<̂�-�o�Q��ILzH�f�3�&�T��{��j:V!�jtfDĈ�3��I ےk�D�M��{w��Q�yPHL�LG�xr=����Y]C�P`����Q�ܫ�� � �B�)߸v%��L�m�֋_��XEZ�D���1;DL�lG������=K��C��'?&�QA�fBa��{I�Eɑ�%�Y%�՗b�~DXu#�>pr Xe�Њ	�|v��̈́�Z3��LD�^��d���iL�v�w�F<��@����,�O�x��:N����B�𖊟(�U���ȗ9;l��E.�����z?5�|����SW��u4 u��Κ@��������D�m����0kP�Z�a�r�O�K��t����z���٨�GuUr*Z0�H.v�$E�dj�|�w��|i������'~�A�ƽ�wvӨV��{,�~��)�Ҟ��I৴|�
����3��$���$dŔƬ�C7H�?0B6�)`�����]q<����y�dN�ñ4by8��ٽ���:Z�3���8��3�ڳi���)C��id"��Hg�2��Ơ�󨮼Eꗣ��zl8(*�`�vX�#1�3��#`�	Lm�Km^�I�=B+p"�b�L�&G��AN�Ӂ������ӳ`�$���|\|�-h��~���f�{BvX\>(�)�����<�o)3�����!#\w�sG��hc�F�ST.;I]�Z�C_6����M_�:�z�n\�ۥ2�4*��ς��?��O��[Z���0�3��l�{�Ϥ3=IǦǆ��a�"Q��^%.�U��I{k���*	L�BdY�7t��nڄ��0?�)�7!ap ٫짿��祃�jY����I/TK68��Tx��w�P�!(�(Q�F1�'�lm&���1yf
+����;0��(�᪝�C�W%��S����m�9C_��?�G@& ����3-9���vm�y��S�<8���E�Z��^��5Wh��;
����wi@q��~0Ӊ������v��y
J��:n�o��}D���1&s�B	ꂀI/(�u�5�����~+g�h��2S-���.�a�kY�f��5��W�T �0|���ǯ4?2���,�c�~/����
|��P��I
Eq�����W���ݦuX�Ğ�0Εr]���J����t�m�أ�[��*XƜ�ۗ��B��'nsC�c*j�=�fM|b�SS\�_�/q�n��R�u�{_��>�6����|e�S�KJsۆ�H�Θ0����JZ6��3Z?n$��GĖ��*�w+�'6hp�i=9��8���Hl���y>�i#|��s[��FWyc���5e��š��5_x�۟U����Vbل%��+,�5�t�?H��n�
���H4��D�/�#�1/���e��Hp��Y��zB��Z�|����Mo*��"%[3a����x����+�-����|[a��v����Ĭ�"���q����	VϢїt�lړ�H�J��K�,�A|ч�i��Qn�=*��P<	��n�݋�]�:�y�`	�IߚD@Y&�5����͆p��nb%��(
(�֕��:< ��H${���vm��� }ŷ&��X�JII�~�
�ېf]DX�2j��
}j�c,��V�|0"��=;T���SJ�@X�� s�r%k�zb�!�d�����囧Eî̧�����H!�k�ɐ�����7�SW��z����w��n���t�� 5������x��B�[�x�1
�KlU���M�u�H���H��R䀴���Z�.Mt4R>�"��Ⓕ�r$��ّy� ��{����$O�J��CxX����`mg��5Dg[�1��9n^�5�gq�3+EU�DbAv
P��majmp'�9M�����`ɨ򰂃u�9��4��6 ���J����m�l U�T<���[�>�c�MIc��T&��!G�1�QV��L��[F�X0?�o�Y�R�ݴ�P��}�x\ߝ-_� ټl����B5�N���Lu���R#h��:`�G����\���؛|P�b�97�|`]%���(�Y���NCm����H�i;�)F�cq'�!#^��Ϫ�a��]�@��5��aM(Xi���P`a$oԒ��ē/���*���ۜ�`��h���50A�gՌ���|����@��٦���11 ���q�D��}W}a����Dy%`�WWII������A|��0�� tT��1t�h�sa���A����/���q��A6�/o�nTX:�g���4�i�V_�픘�ڿ�'����:��H�.o��E��b�C�lt��@��4R��\�(�_�Ϭ�-(��/%�� ��ű�\_�E+�H���� ��X���:��7}E��h�n�N�h�������fLM�Vs�0`݈JV��l�g��˭�k�
U6$nI�J���VQ<��,���Όڸv�6�M�{\�v�Go�҆�(6GxǾ���j�IF~X���c� s?���(D4��7���	=F�?�{p�ե��\hIn�mz��`����)y�	E.�@�Z�%�A�����C�l�t(������Dٰ�.�L����*�#b7&d�<���ً����ϠB�t�p�f�ǫ���A��K�uF�J��b}/.y�_��s]�]L�ϩ[����tW`)�y��K���_!n�N�8��ԕ��ܔSEwzwn�/±i�J��m��d�)e�2����}�)�_��{�qY\x-dk+�2�����G�m�U������\F�����/ �8���#T������ױ�6rl?����l5���z�(��-�M8����:�G!�-�t�|�=�3� ;ŉ��T��+%(l��o�����i�dg�̎7+T!T�ݠ��,z���� >�S��R,_;��xA:�{�;�7��ң�B0w߱�*^��Q [�_u�d���	N���??;�(�4���������h��~?��"h8ޜj �P�0�O�/�Y�I�c:N�ٺ����-xm{�������*�ӭ%0h�]���Hs���/�{���Z��(gK`�
�&��%{$��[R8��H����q�?}�:���ǽ�d�+F!���W}*�x\P�ͬy���U��Z1e��3e��մ,#�W��z�ē���FI�s4�^��YP�	^z �����#~D��}V�q��/���aHUB��s@�� 3�e�Tœ��-봳yrC���cͲΟj�_o�	���k���:C�O�/�H��n_
8~f<	��{ �RN^��PD���(�h(�"�w�ײ�>f3zE��e��`���万0g���O�&/����(�'���T�dSd(�E��@8F��}��(�8-|�������1��R4�&?�� wL��Dp�	�C�Jq�G�4�lc΁�=@�"!��9Q8s1���пjV�ۃ�A	=2�e��A� Btlh�F!A���q@^w��A�4l���o]o`������q�ǜ˅�)z�6�
��v��J����L�x"HyQ=.�}<���F��T��U��R�#Ǧ����X�����z�1>�'1��ؒ2~&m��)$��f'%���J�,�\�}��׶��>���-�x�Z曓�"���79%����}��\~�j͊��y�3D9zܢz�/��[ڲ��;�U~�n�2��k��P"��Q.}��Ug��~d�\��΄�����p��z��a�����4G�H���Rbj�'j��s������1y|iL�P�8�ݪM�I�ME@^ �䌘3IH7�#(پ�`.���;��h�y���o�\FO��#��·�݃����.��:CU��.����㶣�|&��F�_�qJd�k�ɃA�8]��)���'	���X!���~�A��ƅ-t��,��
�]�ʈD�Σi3�a~i,F�nd��}���Ġ��{*�xU�&���8Ej��.�c]$�m3?�FJ\�[{]=Xl�E��"��4����\u��iY���,%|�0�ZB�`������<?ѐ�{!����#��|(�x��-�O�b���ϊWCO�m��e����r!
�P��A9�i�/��ߞqh�^�� incn.��J���j�f(����E鑱X�$@�
?�����W�g�ƛ�z�9��Τ��Xq1_;�K��o���W�h-z-�v��m�׌'�U?�$�rƜ��p�}B\7I��8�<��)��j��H0D	���pS��NtT��%��im��}]z�| ����ʍx�J
���yZJ(|&�^�h�\G�V�����*�?����t�b/!�b�Jy����d;/nܹ_ڱ0���Q�bm2&	�(�a��,�z�8>*K4��-�l�81��Ί��(��Wه� �_��2�G�4
��?�@�>C��$oa��ߍ��E���[�?Q�y%�c��a����~�K=�=v2�{��L�����_C�����~jďV� �x���v�9�����he��J	��?/���l�\ w�����Ľ���C��&�8ԥ4d�^���Nw��{��#�z�G%㡜�S��!�M�p"�.���̘+焊zǳz�#"E$��am�₮��h �Q<�
�{88�ƀ�����%�=�g ���m�4�Ԋ���V�(� Zެ�^�d>^n�An����鄢\�m8*�mن=yoR� i�ZEv�^��;uH��ͧ�E����s�t�L:��3%���r�8�wbM��~�d��CM�n�Mx�m28em�b��o~�;2�vUs��,Y3�*C�.W[H�X�N>q�#��)��E��Csڊ��y�����#�#��8��o&ݰi�!��	��7���0���Pf�r�wʍ�\�����[��VL�s $w䴺���~����2F<3����_n�<�kb���s�lOUM=�꠭~�Z��:�/����_Y��~b����svA[��J�j�����w�\s��tV�B���³�����W�\�2��m�<��"�}C-�� �H����f>���͚"��qe�d�k"~���9<ÿW8��"���db�^��׉�_Qvr�GL��㇔X��2���pf�Fu�q	�^Շ�DBӚ?
Τ��uKB�)yU_�3����hg�b�Lk-VK�Y.��;���$8��<S������gWk����hec(i���Z���0�����"�j�͓3�/�բ��E���Y��۫���{��Y�K�OߌL;�ֽ�H�4��#4Z傈��7�9���� �+�����h�=1��2~��@���}<X�;��7����9�B�)�L��t�-`������e��z�~%T�%�;��J�X~����Q��|�`v��zxk�C����]T_Lt�xc�'lR���������>~�I��܃���@�dN%�R]��}��B����$K�xt��B[��&�90�U &@,���q�i�cC���P+vU.���(��U8��)Mz�!�,&G6�P�쑕�}��O_oZ�(o�"�Hf�� QŎ���/�jJ���[,18��Hڢ�v�qOE�
!^�������Z�#��'�B�8b�� �~��F:�#�);ۮ��h����7�bK�r��_ģ��UQ�01���g�t�É���q��j���-ߢ#`�w�g���Ơ�}3��f�. ��n7:��;%�>1mG_�{k!���:"$��{d���C]i� �lݴԀ[�K�#�tҮ�	�и���	mx6�euK�3�/�Z��b��C])���~5l�����<	2ne��?�/�d���ʰ62�;��(��W�$��~xE{(H�}v������Χxt��)��F���dZy�H�"�r-^�X-�\O�˛]���I��ZFU E���{��o���=��U���QQ#/�$�/*8%����`��,9����i�$�V]\  �=U&;Ñ�H���ל%C��;w����Ro���p�=LB�Ȳ����Zն����Q���_�ǂ�
&��f�[�;��W[��q���D���|��h~Ϣ��b�!��%��\(4A��I.຀�I��K�.����vIػ�+�t��x���5��hx��i�C�q�e��
xR�w�ZE�B�s0�E,��#�&�W�C6���~11J."\������Y\	$�[��Tm��� ���y��C*%�����t���������}O���O�f�B�}63.TF�%1Y
��^a��أ�H�r���RE���V��"����ݦ/�+'�[vm΁�rn���mmsT����ͷqXIJrx�������b+@��A�̉໷�(�K�u�@��`�C�ss9$ �P�
'�U�02~���"����J��,]�f����a��P�R ����� m�´8Nl����]b�7�!
��B���e�RE;(�f�Ya�&_:b}�������u�#:�I:�bV�$]�;�pdzh�"a�G�*��oê�Aes��ɚ�(�fSb��d@�{��i#n�"� ���(�A=������=(rs��`?�+�)���#�]��:ni�p��Z� K��	����I,]n�Zv��Q�J��h;��6����;h�k����AE��(ޯ6z�~��ݟ�8UٶWt��G��6�w:��Jm.�������	%����51�A}iKo���@��[����@�����Ο�+�����S�Zz�� JM�&�/��,ـ��%����>����� m�	x�����Mk����mz�S���6�{r"|� 4i�L�������K�Wݔ�b���c'�%p�8��ꔐ���x �U+�E��Q��A�|#�leh����M����N��X�����R�,��g�7͖v�S2������ &��]=��{(ʍDb"�D)�F~�Q(���l*)�ۻP<})l�x�&M:�� �EtI��GJ'Õn�z�0rH�"�[75;��F�����"�.�Xo �e���j :����H���kbh�cz= ��?�v��nV��3�</�lb�Y&�;��O���p'���N���?���O�[��g�2�KY��q�@c`$���=����E����;�j��ߋ)|�S�/����7]��Qj��P�ft��}�����D����Y����c ��wj#�`�"�8��Ѯ6:�� e�}�{<k9c2"k���d�r�򺊤/Ol����myC�+S�ܚ�����	ßi.�E����B�Ov�O�>�by�_�Cd6����	�-�\�wI�Pa�y!�QlKZ���ߜ����t壩���o��8��o��`��t��n''2 dL�a��g������Q\���o�f�X��YĶ��0*�6���m��3�7�~&�L�і��g֩_� ���Q���B?k�`���kt�V�)�4&IGf�Y����Bu4�+N:��j���b��[n]19O�6�>�7S<4E^R�`N��Ћ���/k�\��gt堤�xEvbG���kU�EN+2���jنy�o1���;:Q���
;F(��=�Y����%�0C����#l�%��K��#C�We	C��#��.ܦ	���V$�kp(�|�R��)��̖o�Ⱦ����Ru���,Z�
�M��ͥ|-�mW5��Ft翑�� %R��o�,8K��1��|����z���'�b�;��)��#|Wժ6>��nE�ñ�C���z������D�k�����u�!��f1܊�@�c���CQ�報��5g�P�+�{�]!y�Cӡ��K뫻-��ot:���n_���C-��w����]���t�o�u7��6I>���֜���"�}�K�G����g=��м]���r`?X��>�͕�`x� Apʆ���"GX��M����D���	�B���0u�-���<�E8��MN�Y�P(���R��8��d#5�I��
b"�N�d �[{o9�4�tO��  LB�qg�]�٢oX���Iv�(L���� ��Q��9����˜E���V�/�~��~Mbר���Qa�%�1ք�1�|��,�K��1���{}�/u�}��#j#��8JB/��j6�����CᠺO1�K~_F����'�p���9cj��H�v��r�'�2��P�<���̒+=z���øgѺ�%��M�Gl8EV�|������u$�����W:@:q���Ȟk
ƿ��%�79s$�jJ����o���O��z$0�2���B�Dؐ�ni�5�`��:���s嶄��,���Y�S=���4d�tD��弾H�Ķ-l��_d�I��F��oT����xn ���������fm=M>�?I�j�Z��y�RC�$~�ޯ+]v��F����2ё&�Ҩ�ܚÄz\?�آ��O�ʌce��w)��k0��m3�������g��v�����|��c�;���&Z�S�Uͪ��]��WD����؟�\1J��������N���t�P�k�1힃0����w�`�b�L�i6e�tkA!�G�C�LW-?�z�}�^:2�M:#�V�(\� �K"Ȏтܗ�.2�B�T�q�:�d��3������k-赬8$��%v7���8�|A���׽\#��i�7����B1���/�����"3,����"�O� �eN�P'E�sQդz]���ƣ�l�6�	��J�习��2�PJ�����O�{���m�8���Fo`���y�e� ꨰp��f�z=F�WG�X�D��-��	��vzj���,���J��?��y�R|pnWs@?�
؉i�{�����aW,�2�+0�ʰ2�I�܉0�qjI	7 �Hs(%�����p!�FmI�1��Kp3	3��IۍU����I:W���
��6������>o|�6̩+Pgx�ƚs)yj�k�s��>�`�Y%"��������HD�F�[5�p�b�mN�0��/�3	�Yӽs	C�;�W�A�*xe��	σ�" 0��@��� >��"66"W��R2���6R^BEo, �e`�Ũs+�lP�:�'���n�;��خ��b�R�t�$
L�ܙ��Q6������Ï�w��M�>0:���\l�U���I��U)>�S���S�
#6��!�|�c޾V���dg�W���*i�]}a}��?���M9B��;�a�d��#
�Ċ5@/F���f�[�rznU� �;c_�{'��V��c�.L��5�Ō���%HEM�ۼ�&Y0��b��o�1J�i%f��^�l9����d�F�C=o��Ş;�U �)نu��|�ӰvXt�~#��M`;z�8~RՍ�h5_�|���}��0�;J������TST  q��4�S)�+��&�&�ܕ	���i���q�k�]��n��)�`�kX�ر�ո���,�B��̛��:��-ǃ��U5���T��s%G�{����� T�ʹ�p�^P��<_p2�*���OɁOP� �2�~������M��1i2�4���>� ��^ۏ��Y+�M�6������$� ʫ����ܢ!D~��9~��|�������v�����>�&D��?�,��|��R��,X<Ħ��39��²�E� �n�$��������ZX��UAQ">�lY���6w_Qg&A�}�?cn�[|Ƒ���4�ڱ#�_ʢ�'/�X��Fn���		3��"z!��Q��a��?7�V ZLZ��h�C�[�� \dx.������h�	q7_bB��Ҳ!��у]9f0��mJ�3�^��<�Lo�^t�`��6�Fr��|�@[����7X1��5�|�>#5��<-؛��?�;O�8 ���� ^4�/,p�,,���(�	��VĨ4��J��C�P��	u}�����O��A�|��6�?�1DN�5����A�#��q�[h|a�3.r}䎈0ҍ%7;r�������֌�Ț�b1�z��y�5���I͕_��߱�B�.�,B� ���(K4�/�^B��pL�@��mEpf�!��@�ت1qVd�I��h�����Y���z%G'2�a�U%`����dÄf�h*]r�I���o�P�2�B>;YmRrN��W�v�okb���%>`w=���6��'B�-c�K�i��s�D]:�p�Np���s��K.�n�6ܴ�F���1y]d�D�Ң����(��Y��y��x�B����`�s�zEp2QC��3�h@������gV��c�/���4�x�]B\� d�?K�Yk�������� "���r��F�6'�_��9-�@�n��f�+�|J����yӧ�:N��Zu)<�kR>d�������S�"�c\⣞rd��:`��>O�o������i0�,��R�z�u�cJQ�D�^��'
XK6�gQ�Nv�b"N
�G7�R[�3s�њ��͟��G�5-�¥�Z	˟�g�`�X��&.a<4
Z��p4s2�Q��=a�j�lq�4���r���B֭����x���Q-]iɆ��C�*f�诎6����P�������$L���W��z�Ivpӷh2�%*��ן�S�A
A�;Ϻ�rĉ�jR.�@����ͳ�����c�%����?2�I��q)�1dOR쾉�A�-��!�ٱ5�(���?�0�J�������DPcW�k#i��`B��)c���Kt"�-ݕ-��[������U�ؿ�L>���zY^�p�����i�pXƎ=��V�Uv�F^w!Z�_��֦����yoՒ7R�	�}����)m���MQ�1��h�%����#b������	^D:`Vm�Ui)*�%Q J^N�k�g����RMֿ�{��W?�A����' z�K�<���W�:�"�㑲bg:}X}o�7"�\��r�T�7�T�P�_�r3�����űpŁ:���J$آgz\�u,�2��@�F�}Ks��nI�H<ni�<o�����oi���t���8�LY��R���^�e�$�F>_�	�xY������8��aA�nFR��LR��m]-�� #U��P��fs�pI[���<��#W���������Y�ӆtuѦG'�[�2��{�m��Z�O�RP��%o�Zדց��m�$�|K�~[�^�ҌR7hft��lY�k��h��꨾2�,c#e]���I��:�e�4]f�D��$�|�:�/r������Q��w���s	��,�a����8 �u�yƴ��B���d ?UM-��b���F<b|
&�zln=K�5���56��c���Q|?@��p�����h������d��Cs.�y��<�O��S�χ����Tz=Ɍ�Y�챲ր���C�)d�65�hs�jh��_Ic3P��WG����I&}G��_ 5��{3� �ΐ�w*q�iqA�u��󍺛#��(����
L6���vS^�8S!�B�ax/�КG��e���*��_�5�Q��(F��ت�M����]8]̦�%cYɱC :�����Ƈ�oپ��fߠ��LZ�
�tc�t�5y #	!�
����迊��].��բ>��~T�b�K��?g�DҌ�*�H�����;^�O��L�o�o�vW�M~ׄ�@)�Z;��c?���b���q��FR��p^0)�	p���VΥ��sCJ9= O��sÉ�,�s���L ��l�OC:���<I��Y9�m���Y�	)�m�5:���[|C�J���ޢai��� ��N�B������X��q'�o�~ 	��x2�7�TW� �����_��9�х[��b��wP����AB��R��(L�$�s����a+M@�u�_���{gT����'۬X^���ZdC1����p�:�<��ʌ�J�GE�k���7]��a����`w"�@�F�e��t��:F�����dn�� FIp5&C6U��S��ӷ/�!ꈀví��@��3�f9it<3AK����=~��(; #�G�+g/�a?���>^�b�V���������@F�HF��|���Ȁ�@a?�D����ʨ��i��h`**B,*�l����3�}�E�&�h� ��+���4S�n�������`�����aضgA�B��ǱP���Ť"$X��h�:qS*�h�8��-u�����wG����?%�it Z��S�v]�$�֨f�J*Y1=D�U�l��O���+�<���I��C�E�z	��tE�h�\F��Vz �w?�c���Fݿ<�p5ס�����fUlOV,���(���E����S� t�Έ��	�����-��H�%��FݡM����Qq1�A�n�گ��f�����<�~�)��`v��JF����ɢ4B�9�O'>d2ed]�@�xDd�;!�0�+���rL��������I>.)�5(��>�8�%d�lMLچ�w��&�g	qK+���u�E�5H�������\k������Q�����M���|)���]�Ä�Bq���*�w�Y��μ�Z��&"�e�@LR��칄��UZ?��)�e���:l]��bn@&o��f�25����"�nd�$�~�J�s�X�lF���޸o��6��HM�%�(o{,F*����?���z����8bAٯ�8Ս7b�a�[�j����/� ������y�ZV��� *��̗!�[�i3# ����0��ڢe�p���fo��T@_sO)���z O=�>9�Ն\�`�m}Pw���Xv�3����D�����j�c����Lkgc�^*������c��� 
��*=&��e��X�:xh�T����ck�cH��jF:�Q�wu=�'RW�`�����=>�2����>5s��f��5F�i'�<�܅Vjt7ʣ���8Ǡך���Ǡ��׈��űz	re�f���t���ch�c2!����7C�>��_��M�G8�u|�}$���ν.���6�,v=��g�!�$C��n��?.��w��w���[j�c�Fs�l��e�_�w����r�'�~�?�E��E�Am����T}���k�Q�C� �p��9�� ��w�(E�fI ��K�6��GbmH┾+L��up�	��,⬉�nA�ƒ�nw��W��I������(ߞ}�5�6O�XШ�aH$|�%���%w/v��&��C��A K3��e	`�E�\�S3u���f�[�p Y<p�l��L���d�R��BY�����<�F��4hI��MTL�]�"���jֿ�XZ����1�Ƞ�e#�~y��!s�۹�t��(7���)����q��U֞�!oHh3�:��������ki�Wb�YU�ax	3Y�k�k̝�B_�/z�}��f܎��;~��,e\�k9O�٧��-���I��~�?tP�c�]nf�g�%��k]׍�Z/H!}���' ~8R�3!���Z��
H~���������;�^���e�`j~��E*���$�.~1���Y0K�Ղ�K2�芓L����npC�	ɉB����h��MRm��3���r�a�tй���kU'k9�*:��\-�T���5,)q������D� \@��<��m�S��l]��������^ L5�&�쵩����R�q����F��(�^�?#G�s�p����+�6k�w>�~���{�eɶ��V�*�Ϩ�wS�v�V�F�N<��ڈ�&`q��U��G��qtOw2ʕ��_%��n���c��vN�`v��&������s��,Mv�JM���d
����qtղLf������`�q@tl%�6�Ӳ����E3t��l<���9�.���>;��!��=S�#�Wi*�PX:�E/WwK�r����GSke�m�r� ]5�r/��jxd��sZ7���u"9��?�f��El�U�K�QQ�^4
m"���(��3�O��1�k����xtu'r�b�,��e��X�Nc�L�Ej��'H��M ��	kU���?,B?�u:@H���섩��3o^ K=b�o,3u�&�	I�UG�g�� �/U��	��l"���Jhι!�C�Sr�����O�i��`��	��Z� 1�UZrrU�>^��+M����?��q]���r��� x��CO�]W����M�����JU�x=Z ��������'���d��<�$g
��X���v��Z��E��ƥ��l���2��J	�OL��_P9l�,Yb'�����mZ�P^����Q֌�Z����*'��LPC��SrP���o��\>D�����i�+� ���/OZr��u�"�K���l�K����|N=>M���\��CC��[Ǎ��.�bx�P����TwA�%,~uR�B%�(������i������ڨz���#���$�O�� �1��c���k��s�_��{����i;�у�3�""&/�T���6_h�jB�V���w�
Q��Nk3�G�1~fP���u츚ګʺ�yo��i0@Ğ0K�H�_>x�h�hrj���S�'�<�4�i�6H�7��Ƞ�2gF��Ut�������x}�|II�ߞ�E���Md��M2n����?c�}���VWٿK�	�����-�#3���r ����65�H"�2�?�pL�k����=;t�C<g�@Z�����TLv����Q�{H>V��g�b�.&*Q~���@Pt� �{W�jQ��^�.i��a��}^���v�e���~
"�f)ǃ���(�.�T�Xo�J�7S����n�li ӯ�W��)3�hk'�/u0�{N��m�1��%�^]3�/?ҿϏ����u%�z�C	��^KR_h[-B�z2���0%�܆�O9�u��er�@�잨����$��ܑ����gG�����zT�`U�쬊R�7(����xd=C��u�w�"�|����O��6H�rV��|$��TlVދ�����o�]1d��~�̜^�EV����Wl%��g�3v
>����R7���1��Cf�V�uB��Y�F��yv�2E�k�[������m̽�>+��꒓?"J4A�5�����F5P��o�r�mi��,��A3�u��y��@;X�2���.�������N�5u���f�CL�g�2�7�Jȫ\���-B����`����Z�ƫ���ԗQ��5��x:�8m?����Ɵs��$$�� �D�A����0ʙ�إ�[�#[�[�9Ѐ��p���"(�?�R�CF����&PR����LIw��F�7��ٳ8��|��}A��G����P��6�/�J�_�S���y�,��,��H�2�Clsڳy�s)U�L�g�B~�lSFq^�t(��g�<SZ��,���-���԰�������@}\U��j�iW>��?T(֏�M��I�l�� ~ �_�&�����ގ���L
؁W�"����X��ͅ4j�z��&��(���I�q��Ö��ɫ��C��.yJ6P�\�k���,���_�	�9��9�g�_+g�	��<�>G7�IN��\(�C\�*ޅ K�.��1�=���-5��V��Se�{�G����}��ԯY2���Dvi�V�n*R�=ʽ�"1.ZR���~�-ٴg��~Oe�s�� ��^"<����>��@����{;��}z���)���i<��Za�����:�9�Aq3��h����שR �k�Af	�.w�i[�h�P_؄`Gt�r�:�?�+Î�2 9]�)Uݚz1.ƚjᵦK��Xc��$tF��G��M"z'\���iL�=R��j�V/o�洝�v����.��a�a�t��a����c�
^�1G[Vװ��)e��pR�oR��Tb�N� �Ac[wY> �9tL���]
)�����fH�o���S����g�Ⱉ`af��#��"���_��Q����<��a�@d���do��\w%7�v@��-'��W�Ŏ�5�+���
�)4NC�Dg.~3��0{-��=z�2�yD�A"�E@�-)�%}�P��:z4b,��{���8���l^�&<�Ɍ�����}�3�qpE�V�g��^`�^���?�$�|*+g�L-��,ߧ��R��w���OB�Qb��=�z��A��q���F��O�L��9�uOG�rPZ�q��Zyh[�%h{�5�g� *�qs1�xdy�:b1�j��+_�:[�M���4a����"T��/�4�*����qs�[�?c �&�]�
�j��i�Vn��>����˶�L�`�S�HŘ�C�q;{�k����/�Ⱥ�e�2��jX5\'��+��Gu�X���VN�Y�ުe�&���|��G������3�A�Y&�(�]`�9q�i����-8�_����@^���e$ ��}{<ck�za��G�01u��);>�+�n	�ʡX��|@/�~���r�q�5�|u�>s���o�H��P��m�����}o�ۃ%��t�煮,��_���.�������s6���n�AT�����1��y׶�u�^�z@T��&sZ�؄�+=2��'�� <��I�׭Dߩ�~X�;�G���$�-��Bqn�X2p�&1���4�oZu��{4|C
�{��D�B���G���.F�E2[S�jݫuZ����VP�7rHY�=*{�{q��e|Ϧ�.~\�t���[D�B�R���{�����L�_YG�XJ{Zo��cBR>�zھ�Ϸ�>r���h��QHB��-q���K%="L�}�"f�%Ei/K�l�*a��*�_��B�L ���T���z*�A����m�x��N@��[�&B�c�?��Kt[x�$Y�j��O^r�vagk�Lo�QoY�$C��EGpW]MJ��Ɇ:�a��A4>��dG���<���Ut�j:��I��kb�)��߉"l&EՏ�~���u�:��m�v}��L�
�k����l��VI����hԆ���V�X�o���Q�-sƩ���������6	K`�e����3F��K��	�����C��8�McQ	~ZRw�lk)�ɗ��UWJ�&�W�	X�rjC���ݪ��Ò�l�M+6�x�s�>O���ـû�l�|9�I�1���w1*)s���;+�u_����[.~�:/�<W;��PL�UF3�~|�@Y�-�@���{3~�(����G�%��Ͽ�H�r�Ԇ6?� ���u|�����g�h?<�E�o��j`��b�M�T���T�|ye0s�׭ ��i\w�0)|�K�'�mܒ_�R���/���	�R�\��#Ѫ	��
ZU��Ö�aꂻ)f���YΜ���f�
XiV�K)��<`�����P����y��嚉 �Y�&�{���e�߭X��h4E�j���(<6A�(d�y�	3���r��ta��R�Evj%��^΄}��Q��@p����Q���k���� ��Xf��CQ�P�E&��������A����cYt#$�j��X���R���(M���_���L�*�9_-��6c�O�T���fa%����?�NS��ޅV/�� �[A�ݱ�Ls.��H���g2�*z�hA�[$�w8����iI_p2Y7@<G�$�к�����k��$!�p�wo-��(�8��@cs��U����r������m�c��o!��� ,�m��Ky�񿳅���.S9W��~���ګ�6F����Z�0S�c8k��?��ʼG
��	N�rD�3j	ܼ�\�Ψ,�����KD��<x����;�
�c `����-[���L/��f�@*��F-���k�a�k��=@6m!�-J��M�jA��d�;�t��#WZ�7�I�׿���j{]���Fo��v��!xe�.(��9�$�'���W�Da��L��äc�A�Cc�j!|"�w��}J�c�R�S��6�[���{߆�މ��F/�)1\C�Ϙ9r��,�ݥ���N ���l�H�����]���@<Y}�?�v�S�V�6)�O���}z]�nk[x�8�1�U?�S�TZ�I?�|LR��1*aVK�ʤ
���=멼�Mw� d[����˙���WY�9�ZJ>@2��/���B@hJ��R�,����T^e߰%����An0�oD�H�+���p$��߲B��{0qK�Wt�F
�:�B��,�)�¹@Q�a���z�dH�	�Ʒ���C�
Uw8�6��P��(1�˩ ~{�-ؘzw�Yd��8h���\���yd��t�y��{^���i�+�U^���~��Q��.����M�����Dٱ�j�M8�����6L�k�k��x��Sz�fl�y��S�f�΢.X��5;��Bk(���ΐ�
�̽�v��dKU؛T����ݏ�y3�b1z6�Ԉߵ��@�U5�l8X��QaI����w�R(�)q׹�Ź
\��m�3 f~���!����%5�Ktި��#pǒ;y�Y�_�,FG��P|����B":��X|#�4�+�q7�)�11�T���n��"��%{���)��^M�$�A8t�o:F��I�0�E-�9xZ���I�� A������8˻vR摒���^R���r��[���
�龕'0W�5J3Q��޶�LF���B�&����y}w������.2�a��nW�Q���� ~Aƕ�3%��v�i,�7���n���遳���uA�O�c��H}R|�������9�i:�Ʃm4������Lg��M"7�|�8�}��.�Db�F-i�&��S}���/*X9�2��w��]��nR��A2>?�ز������t��i�;�c(u�a�6�L��\��^f���8�jo�㒾6�}��,�^��G�`]	uQ3�s���d7`��Q�f,� ��mu'2#�����ԛ&9q�x���>���̯�[|p���W^�7�
�UѴpE�a�#R��Q/a����:�����\v�x{��_GnP��"�J�Cp�����k��J�E�nMbZLN���,i
��o�,۠��?F����6�^4�c΀�d�zU�+ �Z?���!��1	��/����)�˔�I�㛥|�:B�4ɳ;����9F�]&�
lcm��a��	��?�gւB��o��jUV;J����
TvA㒜����G�:����xu��Jx���2�6;�T��O�S��{�#y6�
h2�-�71YՔ�͇���d�Z�6l�#���c�'D���/�S�<r�Ā��'yp�8]�R]�ΟJ��Ҫ���1�=�oV���S����^���T��f<���t�P����_��*�B����؝���M�|9kO�
�������|�Zɠ7?<'�ByH���X��c��(��`��[G�Nu�Iz�~ߛ]}b���P�c$&����hlj\����r�ᖕX�[א �3q=�kv��:u��-꺈`����t��;s�.z��\w����!�7.?\��U8 f���F�3XHm���M�!�@�(̓�&��Y�������UCL^��
lp,p<�HD��|xz�Pq)�	�����wg�����M�m9��ɜ0�Qʴ3�HG���h%hA���[��t_�z$=:���NٌB"��n�����Y�S�U/�'|Oݭ��*A�p�\��`�W���'�l]s#X�VTɯ̓���G�A��J��g��H C4�� X,��GG,x�����ֆ�n ]�5��%���p0g<2���r�M,�Dȑ����u�}#�zƿ�NcOC�����~$R��e��Ț���O�疝Mj�(�f5���`+ !���a��V�Q��[B۵���G3h�/s��:�w0Q��M��Q�M�U��,�#mL��B�5l
	4�8����	e�w��;�_*'띬�qk�'������]�	�I9��A�y� ���/e�<O�D!2ш��'��ٽ�$$�3�7�RK�Fr���6	vנ�6��}��q�T����S��t9֦��W�	���"��^e��C3#�� ���������"{�h[�kw�o5eD���m�fV9P�����[	J�[v4�t"ԋH�8[���o��|�NԢ�������W�<)[�ԓ@�9�L9啘P7LwCȓ���=M{W�x��щJ�0q��~�WCf���f��of@�8��a9��zar%v����ILm0�.Ktw��B=e�by�MI4��o��q�����x|�.�J�L�ubG��71�D�kn�h7i�Nr��"���r�:(��?D&Lb�||��B�Fh�1 #������/Oߞ>�k�O�DЦ:`b�f�2�"kt�+��[��äN;��p�"�T&��^K���̓y��,)�^ԔK��>����g��d�����;ٷЪ����¶Lެ����Et~�'�d1�Mv�˳�@������;c~O�l����Os}~�V���n�)���.I��b�I�G��X<����G�	z!��v���u-dR1F,���J1����-���Ĺ��w5�iRBh���!��_���a�B3��4�����*��*�k M����"Q랫SSEH~��܏=|�����|��ڱ/ Z���	c����JS�q�����td��Y �����H�R(��f�F{KE��;��S��{�?
�%G�d�z��i������(���^�����uI:�:ЍSa��q��x�"���� ���l�R�7�'_���t�H&�Z����7m�aD�f7�e&�_�}¥\=3��^a񤕵�����~@ȎƗ�[On��9c?�y"��˵�rTѱ���)S�+܇΢⥶w�f�£������"A�q��������X����k^FY�4���zw�7�4�PH����ڨ���D�}8h̿H���^��]���]�\�3��Ľ���MO��c��?���/��5k`��c+3Ϋ��?�3�2lp�#�x����ݢ�n��;v�U��<���dE�-���� e�U#�ҭ���a�'���G�#����'o⣀�8$?�@B�����֦����K��k�'�F� �8���>��t��O�\م_s��ni4��s/R��y�d�Ɔ�۰d�ݭ�k	S㶣.�yY�}�0G��QW*��1$�~	8	6�!ؕ�
��29K���6r� ���~qi3Dsj6��H�;+��	��.���q��������F��񀜳��!bɱl�ۇ��	���˽WU�дϫ�>������9�3�O^j��*��������oF��z��nFn�p�ƛ��#]B�o�nIe���)�E5�A��FjBk�F��9Q hvMc���}6d减Ǖ�0��A��D#)怢}p`7����������5��28k�᢫r�Fԯ�d*pl��#bf��Ii�U�?a�A<7֛~>Z���=<�}*���i_����P"0��h
4�*�o3�����c{x�6��E���bBLa�1�6��r��i������?=i- ��n��Bg���9xʾ���{cp7>����Z��A��R�[�	������	tl2�Џ6	�<����u�K��f�̕؊B=׋8�hC�y:S�%v%��-�c�2���P�K��?$ASz���w
�
6��ޠ蔣 ��:T�f���%h���x��ő��R�Tk|��xE��52����O� p'�n�Ð�Y ��F�-�����E�U����x�+W��6 �2�@��& ��}g��\�}Ǖy%��mqW���L�G�n�ܼh6`Sj���R�.
ss���4�m������J�xA���)]���鐿M�_�Nn+<�!�5:Wooy�_H��H�U�9��h��C�6mp������5��Q}�$���rq+c�\�]�vt@��h���5o���Ȭ-E�s���Ip�q�#�=i`�:n�Gh�#�&��i����}L��_2Mh%]-�X5�j���������z�Ƿ���R_�&f )�\v�O
�wOb�!�X8V�N�H(c�A��F�u(T	Z-�OɅ��X5XX���䷆.ש>@�*��%%�����3��/��U2�-S���(� ��ݳ����|���W'w��Zػp��bu��W�>�,u�\�?�M튈�ϝ����=���b��ܢa3��C�#VŏФ�>�m+��Z'c���(!�'��j���(��u&nA�}�:3kG~w_O�7\ѿ��!�K�;�MLKo�������>'���Ҫl���'�$&���P3QG��U/���	=W��x�X�a�������6L�� +G`9j�'�pq�?t�pg���}���I��/���2�+t�wH����%�K��S���7��OCX%���t� жz?JkM|ܺt]���ĸ"��(�/�y���xz�`�K�}�����xX�R�ga�{����⏗;���zf����/M�^F�!��=��0�ltMXo���܃�#��<p,<��� cK&ю �[i?�������å
���2.$n	���|��h����c1|��b�5�����7�?���ٻ7E>�M���/5D묅��~�u=�۹vJ눝$I�we���_Ae(���Wgj]+𧬴&��^�.r�H4	3槐ZG^��� +�gF�#W����C�c�����C^W
�Qt��y�Ƙ㮷�����{Ʌ���7LƢ�~������j&�L�c,�4N��,0Cҵ���٠e����%+���ޮ���j�v�9(���x�Q,��jn��0y)�
�����������%�"3�&��!�v:��9`�R	h<J�/������֩�W�q��ה�!g�fJ�
�-X���d�a`6�����]�@̤:�ϕۉ;��|߶������h���VR���8.�SF\QS?���4�}�3���,��PD�1���Gwݱ�e!%Ϡ��B�Q���?f+�Z:�
����D:ˊ�#0M�X��� �!&�<KնB�Ģ3x�
),�����3:M�j�=�
�����ߪGȑ�(�.S�1�Γ�+^)�N �$w�Π����6]hl����t���4��@$��sU��\_sk琠�i�.B��*��؍4�V 3>A_�?�����Z�TD�m�7H���L�gZ���d�	�`��ɿK��2v�!�#��pU�X?��[�i�9�[��ga�6��
�>�c�q�0~֞>�-���H�Q��	6Lz]e�CF���?�]Cy�u�}z��D�E�Ĉ[=��������T4����/v�F�oM�"��Cdp���3@�������b�旎�k���AϘ��G��Y�7ByxמER�d�k|��~.�L��w��{Ez�.q�MD�G�ƁSuR�q��XM�������^�c��`J����)���6�S�*	�G$���נlw�F�l�����gTͻw/��rV6n�"�Z:�l��t!��}��-�Gz���^�)؃��� � ���Ҩ�2<�\BO��Ũ�kB�f�
Ir��r8Lu�^Q�u���1��:�c6�`��	-Ro§�5a�ƽ�߮[}�j��eC�S�S��&e��I.ü&�����!X	�8�<Y [:��p���QM|�����UGC:�
x��ͼ�`�<���t7�yu��[}���[�{a�_��?0��Dc����w'�H췎Ѥ3F�˼��� �cJ����4/��u� �oN��i�
X5e�0�oMI&]r5�zvUn n��q$���������Ky	o�՛@Ԋ"��� F�����wQ�(E�P��,�������&aV�4p�W��ǰx����(�Ar�uh�	�X�����F��m�}��}�̈�v��r7ޯT0t��X.{�S*��m����Q��}ު����D%�`6�"����ܪitU�͇��m�XF.�Î@|Հa��y�1�q�\�l��싛��?7�!���bc����{]ʜ¼��*FŃ�q��<㮮�Rβjkՙ��â��%��L�M8f��w^o�u��QC>k����������aW>���c,�Ǧ�}���,1xAñ�8F�F�֟æL[E����qOX��g�]z0��5�*���!�×h��Ko������jS������.O�U�N�;�:�V�TQ6�Fbг.�$f$�����_� y�)0�qj�;T���~��K���X��K�)�H��9�=Z����	�J9�㊶�R�(��$͘�e��r���>�' N��4Zcc��R-G��io����iV�zbU���)��is�6!:�C��t"�j)c��T�_J������Tq�ۈR�X���4k��:���S�z���?q�!f U��wq�u���Nv[L�	1�XA]P�݇�#d�W�l_���[_���=ߘ<,���tљ�|s��%��]��R�;�y�r;�F�|t:D�� ��n91��E��7b���wpZ��ס�O�e�/pd�;^��k���:<L�/��
���v�;���Z%EsB�
+�4���ы�E�ۧں�$=�UyC�-S:�����u����E���Ӓ�pU9�QqBJ'A�����������UX����`��VS%�x����Q�3_f^�	R�u���_;pI����p����X�?��0�E5Z�"-�Ք�D�E
���k�ӷ��T��kѠ�T�)�� x@d����`9�������3�јv��d�]�O\����3�O�F��s�MnYq�1A�C��l�C�����[v/��y���u�����"�%�~D*g��}�Rֈ0�`е"F����������a?��b�P��%���q�X���xh~���6�b���7w��ogr(����Ox�.T��^�S2��t�2�p�`��*�RR>�Ƽ1�O�_<of�!���������,z��YNTz�����iG|U�����5-��N�Ŷ�+#�+�pX���� Jط^��W7u75��l0�^��#��U �,��W~7�rg���DYs�#ys�}� �����o����h^�b�r�8,�U��t"|�Vɞ���r��_f��]�.�k�?�ox�촑�Ob_���^~��dw���"�N-��'�L����|�A��G�o]��*�6�nd֫��c:��˓��y��{w�$��l}�[Y%��L�6�&�<4�=3kZ<!�/yAH�-9����
�Č���!�	�5)y�H�y6>��M0�m%�A~��z���S��k
��K��5(��E�LX�'�y�����hӸr<����jm����v��o�V�#��}�h��yq�/��E�����݊2��w�G�|q����	�u^f�\{�e�H�.���N��1�H��T?���21I����`�M������W�� q;,V�a�B���wV�1Ң��k�W�W[Ǥ�)�na�7�� *�q>�ժ��&��]��T�x���p:<GI���]�4k��:Al���R�Y��/��l�b����*7t����]UZ}��	D�B�+<��&�3K-9�
7(����zm����>�2�ol�g'�A2�*u;n3Q!�؟��y���.���kő������'�[Z�5�#iξ����By�%���w-���
�قL�f�9w|�X���R;R?<1 !���4A��j�J�z���	E���jcbȬ�WS�e��|>��5ѕm��;��٭�r��_���i��d�Q0��z��Xu���`i2:v�Ă���.�6��\�I����b�Gfq$L��E�14\o�qb�'�с�:�s��T�$��Zw3�d�Tj�ꖨ&z�p�<���.���kΟ)��l��w�3�d�d��J6ެ3_�P���3���\ҟ�W�.JT�q(vn���@�՛a�|�?o��@��D�� ��J��Y�ʰMZ���֬\�Ym6p������9<���-��1���1@&t�Z�1c<��r}�����Ɇ|++a�[��(_�x;cs&��<��e��Y���:�֙��8�ެU�&�<���Kx2d�� �v��������)�0Xm���ƫg��q����^�Z��fN�F��t��<��S�p����ŧ���򃻣s�ق:%�j��B�����xK�\�R��h��&��u8)?�<���:���9�;�'�����H��t�f���3�s{��ެ����g�FP�#$��YÕ̉𘭘�Kޖt��J0f1��O�f��v�"u��nyܝ��@����K�~j\�3^�B��@Ґb$=��`��n��eI�h���2��\��u�K|3��U'7c7�ѱ�����&W����Nh�sT�����̦������r�('4Z5���^;�_�@U���qz�1Xut���ng��_�tp�Cx
�G�a[rc��J����n�����x��_ϟ��]�_e�jyU�2ݪ� /��Z.�j_9�uJ���?lT�<j�U������O��YXW�Qg�_�h��hc�i+��ƥ	���&��L���}z���d��G�e�FxW��������*��PEA�?�ߤU<�{0$sT
o~�YÚ��x��l�-r�%9R��g@
�R�p�(Q(��E����Cof��{zF�Z�e�L]��
�� x���@���7HaBXI2m����f�_���� ��PH9��v�(� �-�Qo5�z(�e�;M*R�$���N�֯�݂����*�CTÌ���(�� ,��,��nv[�q�^$w2�]�§Т`Ķ�,J��茥M��_����aҬE�ZJ4?���8��q����.�h���~U��d(�{�!q��xR;���k���'�f�bV}�Xo,��5(�ʉM&�4���/Uzc��G����F~��,�q�mo|�����I+���]ވU8+�q@� ��CK�a��C�6�K�W�aK�-̴�`M�ꌒ�lN語]�@G	�@���SJ-��z�3T�gUe�|���%Ҳ�k��p�6�/��4]�6��R�<1������j��T���	�]D�77�"������Iw6�?⬝��ମ�ֶH���d/��|���ԍc�;��m� ��Dq��k��8RY�>Ҵ6�Y"�M
�s�ZE�G�7��=I$]^����Д��m���I"Q}�ڡ;0.6���`q�U �A'/��3't�"�"#�	B���u 	;��E�m�r�Љ:��=����X/Iby�̅�{ߔ�d�mYyz��^�w	���hG�&k��F��a����`�*K����U��<Z��9�v�i��Q$r��K�8Bc�����! ��O��uw�Lꋿ<���Ǆi�v� s��~v�:���z���k��3���;�wx1�ѲGu�^8�CT<;.��4���Ҽ���R+��hJ`b皥;ț��}�.��}b��} �M_��T�z�,�S胣��n����2��Z3�����H���U���[r�`~*{k�H���P��*oCn\,"+�8��g�޲ �K&�ȯT�b���l� ��U����#^"M�B��-�%<W���@X��zB�p����G�K�L��{43kbH�g@��f�Tb�mb�
L0�~�n����_��Cc���2�#��ߡX���,i�r��G"%�5s�A�9�(^@�� 򙌌�^'vZjk�lC`G�=��L�1��PBc6�b�W�)��Ρv�&��C��}y\ 9��h������F�(  �,-�P����̿w	H:ԡ�ԕ���d�i#5�&~�M7~.4$����J������Xz#��qh�������ܭS��ad�S��v�aQa��V��*���ci����G�m�{�W���G�4*T��Vw`{��Fp�j�{|��e���}�HS=,�U�����:b�Kn2ң�q��]mF'XNGT��4J�����c�=��/��N:�/�f}z���(�9�Ă[0	�~�V�O���Vqݲj=��mj����}W��� ��`~�K*�/Tr�'#Bs�Y)�-�x�`,�:�D��*�ni��G����-��(|%%p���N�������H1�'�J��)�	�A�^�Mr��Ǳ#�}3��_��c���Y*�8�= F�y��Uԡ0ˈY��O��@�yxc�����&_2+iׂ�DQ��˩����q���b���k�!\���H�og��b�e+�TH1��,�F^*椅��FA�K"J[b8bD�<o�	lm�﹈�z�����4�m#,B��#h=�������L��kg-�T����R�a�x�J��U}wd'0�mzw�HU~��@��!uë�����SF���҉h�vپ]@y�r'�#[�Wli�XO�w��o|_����iy�*;rP�p�渰HT�����7�h|��)��6�F��J�����v�tT&R�^�VǶɴf�,��ǻ�``�1��`CAnkrL�w���[��Y�����B���c'���Fj���HED��2< ��t�@%�oJL�軋�߁�ʁ�4�f O���E�ba�D�׌�2�RiEfޘ+�l&�xڽ����G\�TMK/��j�	
×�?�h��Y"�Y`�̟����Jѕ��5_y�ym�:m]:�R��p(툽M��9?���Da��W�KȒ�<�V,L���k!����g	!6
���vF?P���vg\�X�Ye�P4h��рB�ܧ|v͜���+<�AU����þ2�M۳��R���y䧮�(c=c�V�0=OX��gїRs���X��,��^E��mf�aCdaE��kbH���DKKdU$�t��=� 4��~���T�d,�MG�ꂀP����9kߙ!�H��`]49'XS'@^��'4���>V&�$�tQhaJӆ�8\��.�c�����D� ���z�/���AuC�L��`��h>px𫁧�n�D�-�{yԱ�j0��3��1�&dk�%o�i@gO �	�?'��2�1x�|>)n��}�oO�������� �0G��V�AEA��/�uE���6oUyW��$P�݁?c1챘����v�$ۼF�>�10����������7��e,-����il仓�E%��^��W9Nrӳ��ik�v�����>��n7���l�$�x�'ȷ��T/����$����Kr�7"��j�5�Y�P[M��F��u��|�hS�7��(���gǛ|9�H<|H�<�g���K���R���bY�N�V<C,���CNifa&�!�x{��.{��x'ԗ������F���]T��k�,��6FI�Ͷ��R�V+#\"�{ ��$�Dx�n
��i���*���c&T�.F�s��R��ԘVW�E#H;ws'��'(����8#$�g�w�
eRd� ��='�R����H���K|Ք9�
�}UrҖ��,T��|�f�v�d_m7�d��/()UR�ѐ0����[�?�s�nB�`I�T[~�sM��B���f������n��n�"=�~���]��Sں�˕���D��0�+a�ϭǞ��K� }���p堲R'��oI��K�U�bmWrr�f+S�`��It�

�i���YO�?MPA��l���'�l�^����)�=8-�y�x��?��qP>���/�*�Q$#\-�f��U;��Q����Lo�)�,� ��L�v�	[�
h� �P9���+��j�ԛ���=n�p�p�ɗɅ�s5
�e�~�=��_��Zy��
�"��d��i��R��dmͲ�n�t�y.��:)�ۥ��=��(�����.�1��_|�]ϋYrˁ��_<�TW�Ë�Sf��c�<Wv��X({l۫�⾸�,f�5�����Q�.x���ֻ�=0����3��V��^�="X[.�p���D��A�t��`�4J����p���{���J�<���j��T}#��*��\A}�ڝ�C^�?�B2�e#?�/��P��	�$�u��e��EX\�J�X,��l� p���'��w;�!*kbZ�En0�8�Q�X�?��w�֯b��Q�YS�|��們����Gcm��h���	{�ب����K��A���#������2pj���J't�˩�f�9)I��y��y%��-YL��M���s=�S"m�K5�m�$��Դj0�ٳ�ތы��uY�5�X�2����;�T�!l��@�a`}�,�aUx���z.�p+��^Og����M2�p�)K���:g ���S]�U�" 0oIG��j�iԆX/�A��*u�>�C�4�$@� �s)xH�� ��tȲ��0a�gtl���h�^�6�`EF�HZ����\p�^�g8#���ks�\���"n�5`(o���� c�nL����4��1�*���ot&�s��j�1K��ƬI��T'�>��g��l;���ń��͵��_GN��9"�Zf'T#1�gho�)Q�Z{��| W@�Fͤ���$JՅ���z�!0�Df���:�#��ύV�KGy%.�K�X���ā�\A{}�K�A�V͎q��(Ƶ�S��Ϥ�Qj�r�Ͳ��Ldإ�y��rJ�T#n�������~i-��))�)�0��-��f7:���
i%�-H~���Ѷ�K�Xa1���"B.9ܕK��*G�-s�,�t
��o�� ������eaaX#d��Ȭ�o
ۑ�<����r, 5/��j������_!^���)�3�Ia�L�k ���v��%�o��I�vF�!ۤ����Ѕ�x�"�2�K0Am,�����Nm:u��}�����*��WC\��$��BM���̐��.U�l��Z�V� ��Z��m O�V��ǖ�GW��i˹�4Is�����d&}���<.��l��XZ��[V�Wio���U���j��p-�Ұ�4����H����!�<�|�x;��K�a�e�� x�gE
L�KW9������8ge��}�HO ��B����0(���9�m�iCן͔h�#�Q�6���2�0� Rjv��.���/UZ�\e�����{�� �(	��ե�Dge�$L:!�@X���^�K";5�Y�O�Y8/����ʣM���l����R�N��Z腚B�ϰH���Ol��h���w���F�r�/,�V}�U<m��3:�w�*xi�����N��GM� �<U�L�����M%�K'�vJ���BFb۫?j��&���F�%'��bGm8v���w\��6�ݗh��xK��Nq|��z�Dw��3�����V��(�,��:�"�}���#v	�2�a��[����s�~�X)�V�[q��ڱ��Q�l���a��ƪU�C5ȩ8��[��G&��^����f��/�����	d�2�7@��>��m��]Q~~ gz/긳�e��}�~�]N���L��V4SnR�!K� �>��͠7W̦��n(���~^��X�����;K�a7sg�)�����5v_u�@>4��V�Ƅٖ��]1���~Q�x�I��ϡ����;ۣ׬Ķ,�m�8S�\Az����A�&�ϪD_�����|�n��f�W?�0����V>��ٽ�*�ƨ'�{~?$[1����H�c�YY�;����D[2N	*�\*��88�۝ۍ�����k��� E��ˍ9B�����A��fl��o1�bS>��+?j������?;��K<�8H�(���^��jy
�`'Ҁ�	�5������N~s8l�����\+���{
��e�U%v�w+f���	�E��ehp�3��w���Y�`�ݙ��LCc�����2D'=���p�P?`�^[�X�<��zG��Cd�ǣM�I���geB5���'�oX�z0	%�hL�������H������n�?�?vy�ԡU�|� �ڤ}��L��nO�?���<3<��SG0�eM�+m�$E�S�E�1� ت�f?X>$O�kY!��'$�yh�r�QV�q��ʀF�\�g��4�Iđ��-ݛ��/~	{y$�/��?�a.Zj ����?&r.���ہ<	������O��]$����2[`���V�
r٢L3m=���;��5�2�f``B@�y~j�H>�V>����M �HݎA-0�q�~#�ޱ���)5狹c�6F���<T"_�>����Oj�o�#�����%w�N�1DHq���g�m_�[�Wy7�͍U�\��U&�S��S����8qQ��4S�#jY�S2F�-���YG�t��F�$������+�r�'�2W�{��M6���B�`��m��	��~�'~�ϖ�B�y����5�F�C��*��V�Nc�[��+/�[h��;nY�����{!�SEOqg�������L�U����f��r��f�b��&�� "̝ٓ#���0�\"�g��I������[&�����[ƕ�	����2���}������j$��4�����57�i=�ۏ)�� �f^[o���40���������쬏z5���K��1�h/���k4������cF�z�9V�#�H����n�1�+DL��}�^��M>a�� t���9S��u�`X��>y2�O���Th�����F�� ��90�i�)�$����Z�S(c�qk�؈�	���5d�9`�|�1&a�l����#$��(Qo�tdN%/@��$s(��y##��5���V���%�z�Qۨ�NK�M��W�6+2�f�D1�K4�i��R`��Y�HH�W�\/!VUEo��乪8L�\>-�Calxm�;!��y]:�zbNG�=_�s��Mu��2*n�;ѵY8b�˕I֯�@��+ݫ	��}g�}Îꛠ�� /m���#���:º�Y�Sp7ż��9`<!������&
�N�ϧS��U	8Q\��#̂5E�0���Caܦ=1�b�C���ԇp�0�,ٟF��r�Z�Cvr�|��>ø��M���
�x�Mkan�#�3��'`B_ R/���W�-�����M��Q���.�g�P��ְ�F��Ƿ���d�ov�dFG�F�6�� �oQ_����A� ��>���[���q�樜д��*]�0uѱDi�9�&̼ٞ��+NF�M�0��{i_��g�_E_
�k�e�[K����!g�`pd�3�X��"ʾJSO]�Ԯǆ5N���ޤz6�=_e�fm��8ƹ�W��� g"��I]A�:B8�8o�b
krq�M@KY�ǟ������Hj�h3zD����QHת�"3��<!�j�ψ}���8���������̱�JX�zk�����lE�A~؈߇���\d����]tD��=I�����G3�E��i=:��s_t�s��{Y*	5�*��wU�Ք���N[$�b�%+���`��|%��@�u����g�A��8�/��b!��W��5�7�w�V�������-�^����.�<�2�{=��1A9g����,�s�yt33t�x2Iơy<�@�ǇR���T�h*k4<�u�!�A�̊�C�!K[���"G��J���Μ'�U̟�C哺��l8��&�P�4P�X�{oƍ$6,wӜ1�Q��4UJ��x�4֣y�V�&�� �8����e���9eC���J?�!-K�`�
�����B�
z�� ��j�"z_���*�.�[�,�5���<��\݁Lݒϡ�p��?����%?���#�#pJ/e>���B�p�8,�"4��$��k�UI�v�xm�4����}�S�q���&�Q��{��k�52�#u������h[h�=��	nc���\�ԯA59���ԫ���T���#t<>��H�ɓֹ�4� �Xu�Wh@a������&�ߘ�#�<a3!$X�H,��\���� 吝�o!W�ه�$���C�C�P&w�v�3X(]�R�Ķ%U�h<�����t��j7��k~��:��笽�UJ�;�� 52�hA��V�G-|�Ț�+�S<c�.�O�ժ7��u�7��t_��o��2/��o� �x�,�֪��݌s�F���5�yO,>����=s/��7���3]8<���~�?�v)ҩ���p�N��º-���n��@/��
�K[toEҧ�8�-o�0f'�"�k��(;��h�iۊ��)�5���������Ad�FD�\6�ߡ�ߠ����9�H�K+#�p����O�S�:�4�iV�᧙st9IS؅"�2�����l	u�8%�����G=VA�D�G%EH�o� J���
�ڌ���R>����c-�k]p�U9`:x]K�ZǛ��Js�ֺB+�l��D���m�E�l��?�h������t��RW��k�6#=��A��Jt�90}������-�O�%�fН�Hu�
�d�i_B��r'n��v�N����P�t����Rt$��t��5�Ҵp|��z�8c�\w����=�|9V����Z]��
%���V�L:�p�Ţk}���2`� �-�1t}E �ψ$ߢ?u����F�����Λ�߹�җm��t�~�q�[��^��ݥ���Ae �:��dqa�I`#Bc�W9�a,�]�~��"���ս�2�p���)t�f�5�S�SjNd�#��tx)^4�{��.x��l�21���r������]0�e�WL�VɽAm` q'u�E{��S��d˘�w4��I����a�1��1w|��:��7x��r�o�tc�!8�\�kGA7*>�KM���b�#�<?���c��<�uP�r�Ved�n ��y��P|� Өn��Z��u��\��<�2q�64�����-��kg1�����&�>�ʦ7!]�ڈj��i8r��O�� ?;142�;�1E/v��>;a�(�7+ !ؓf���82;ȹ�T������~@��%�\9-���
�b~��լ^�X#�WU��^g��{�|�����5G}��w,2��"G���
w<y����J��1�L� �n�hs�c
���� d�]T�Ӧ����-�֟�Ͷ�a,�EsZ����YC�0?�G�:Kab�rFm�9dJe�i�$=�a��njvv��h�@�atS��7�W�ץa��J>9�}A�R�����
pJ$n�74��0- ��7�����XD���^�;#��ƥ�g�MpYXd����9z0���uA�����=�[%��k� gf�y�V񧮤��w��4�#w�����`[��+o-�mL�oi���:bkHy1�e��I�B1?��B|f�+�����V��%Xצ��CPgG�!�%DM��`����#�Nx~�	A"�5ؓ��@vfx�.6DJ���@e�ءU5�������Ɓ�Ϯ��.���9��2�l��7P<Z��(��B%ܴ����E@0v������=�rոB�\�-Ўͮ�h���WW�gw���7�����4�B�s���+�=��ŦV�I���l�xF�i��`[�����ٳྨ�N�$I_H���*���K���]��]����rc�V����1 {�`~§�D3�5��d�[�;A�p���9-d��l��AieTjDU"��cPR?8���Lq�����V�׼-�I���oʷކĥ�4+<~�<����L�~�I�u������-�W��k�E�Ť/�X,����fp���β��A �	x>�J�>k�Ėey�&������̸F1��ih��a��#� f�Fz6B�����%��;;�`�
���F��n-ו�"j�d&��������L���q����=>�A��S��R�2�pj;�?�η�T��oAձ�=\�"BQId����\α��\�����)�{���~�/�c�SJ+4��<Ꜫ�B9ޖ�X��É�x��I�f(a��@~J��Ɣ��~`B�{;�� ��fh[/k,O��������|�k�y^�*�6~x_J:R��E�34B�e�V�����Z��)\�P�|Y�T����YJu3t7w�������J�t����t]�9���p8��V�Д1���e(S�*FW���gL$Tx_���RXUm��}(�@j�C2ؠ�tMY��\��cVX���=���[�qFl��"R�Ǽ��2�>���J�5ܗY�JX�k���]uh��z�Z�i\<dx�@5a�$iW5g^�_��`��U�Q\��kD�����
^�'����d5��
�wuJ�q_|"D?��og��PXY��������U��A�ٚ���?{�o�cl�$��=�3�sUē�+dL���=����s�&�w�;�pnP�#���H��Tr�G��х���n�r`���6#�,n�����J۳����Z+�#�M�μ_�H�]���=+d��v<5I�6)?:[ ��n8@�d��ƾ�T��M�t0|L\��M��?/3���wvߡ�I~:2ݝbe.c%�K�{R6�`����<na�8�,���%����>��2�$���M�=B���,�� �O�y7Nw����VA�4K8��h�������s.��ˡ+]�"�Y%L�m	{�s�R� �RDluh7��S^�>$���싫��>�����ԡ�VjD�����AM��\�&~�O��_�^=m���}�4�0)
���1p�	��r�7K_B&?݄*�	�J�T�*���g��WC�n�`r�0v�>4��1��o2J���p�H�Ҙ����7+�2?JQ_B(!�8CD�u�a�ݏ *a�����ri݄-u�S���p�0Y�����9��p ���[�>�O���%=I�qcۜ�,M5_a��W�\٢�X�
j�Sm~�\�1uѰa�F���X|��~eq�D|?�~�+��`j+�u[<�Z�-8��M���8~�t���)�552z�u�O�[���c�(�@� �=R�Vr�n��pjre��V���=�x^x�>}�/ڔ��ȿ9%4��I��@���׽�s}T[�9n�jF����|:0,L�Ьuv����*��������lbЁ��BI���+�|�2�>���u,�~F���$s��C4yN�wֹ��$M��2��a�s$U�߫�Oo�U_�����&n�5��E'?��H_8z�߿2�p��Tv[\ѣ�7h�;��yR�P>�_/��w���-|ʹ�$����x�A�Z�*'ĳ91{wx�ٴ��.�VX��̪1kh�1N���J�.�z�TrZ��TT�x���3c@l���.����<�H 0�ۿxG��#v��e�>}�7�0�V!1���V3��;0��4�f_���赡#�=˒t?>Z��fBҍ�.H$���.�4���WQ��9�"˅�=�T���{1�-B��h
���g�JGf�F}��":�(�P��~Z�WD��M�%�m#�(Q]�s[v z���% 3ߧr���Q�پ�9�UA�m��mm�FhUͺ �/����KPk&�q}������ٞ'�ϕ�[ɇ��mݗ~�3�����j4�V2�)�I�&��NM�8��Q����m���GVp�>d,��w�l|Lt���nߋe� w2��<|HbK �����N�1A�m��Y�-�F����뀯?���֌�?L�$òN�گtn�B�n^�,�_U�3Ƀ*��OV�pjEŅ���NMQe���p�9��//�\(�Ь~:[*���G�X������$���>�iT�mC���î>�^r��U��x�_ �Z"�c$2���3�o0�O'��ǜuz��S��o+Md��� ٖ��:��h�.C��N�&�ʂ;�앺������Z��mB�RU/:0�J��0A�35� ��)��t�m?D0��`\1�Q�����,Bj�Fk#���J:���d�U-١���$�	� \L�oUN�z�k`Qa�\��߭��M�6#�ߚ�����k���������X�x�-=�Jj��k�������i�ωE]Mb=�2g�&0��h�� pȮ���r��̅�ș���,�NV/�KT�Ȭ��T�ĺ ��3"���ryAk(��k��2���L	���:���g��(�e�H}U�quم􈭢z�%Q2�`ڠE�~$���@���G%��Wy��jGOf�D@#��
�#�֓�3�s���R�_��Li'C��K�>[;�^&�)E�~0Z�9�H��:v�#�޸���K�+��8��Ӛ:��W��F��nUF����9�31➜�/T�6N޽޹�������PsP����]��U�	j�,���y]�8�� g�+��#<z1�˩��!�c���o1��R,���@��'�8�M$\kNU��5〚�fV�ӾS���_�KL���D)VDN")ħ�\��g&��� /T��o8����{�gzPQT�%%�gMB[3���,*�����x
��<]�6	.v�0�sWluO�(�&`]����B e���Ȧ��^��.��:��U-tF�K ^��o!_���8(lvx��*T�0!?$#�/���>���;Oث Q�غP �Ö��#{��}`�K��[�0��`B蛒�R(���J�5�ķ��'�ڤ��0$�?y����1�3�pm���Y���[�@Q�B�+�qߥ���U��5z���,pC�9���}DeNaɂץ#��TX���jP�I9����ٳ��p�%M��qt�}1��X���!�Jju�Z��v����}pt�-x5�x#	� �#;�W��.D�[�u��bthf�Vpں�FI�DS�c]�E��P��m�ܘҸ�	�8�1���d+9��ۋ'~z�>�Ȩ�(!�6{��)�0�
A��)5 k�
�n�\G�S���m}>��[(	�<nB���6ކr4�9�\L�ޥJ�#�I���a�E͘�q��Z�0���?M��{���q=:�P����(1ȭ�w���x����x�����1V�b4��LL���?Iۼ��H��̬}�]&����u�l%�����>�J����S�8��<G�w�)5�ԫ[��Lީ���B	¢T,�O��B�o��3�[�4��W��ɤ�Q� �$J���9���-׀L�Xx<��KR�\�7��y5I}�1�}W��N�l7�b�#�=��@����D>6RY�z9Z��~W�J�e$�!���#,*xn�I� v�k�8<ڙ6OO[�vAxG���Y�5eȌ+І�Jo�w���)XL�	�c�����3��/��:g����׸wO�G^U�V��Q�������p�M�5�f��_�K�R�.�yfs
��$܌R`�f�$�EU����[��-�G��'��Xl8���T��w߫IA�򸓘�`��[�_���i�B*s��##@��^�Xf�n���|��:���[X��ϝ��Mk�����b5��Y1�j��yrZۤ�;G���8�_�!�Ҍ9c�&��h�,є��Y���QL���G6F�gI�h0vS<C�V��T1/2�t&MH�q~E̜x|�(q+'<a�l����^�N[b��PNeJ��O)	U�,�A�0�먾�$�U����>���(�x��A{��(�n�l�?0�0��!_'�8�-5A�ٻ�,}��5Ҝ��h�����L0��,r��s�i�M�_F��@�Y�1� 1�@��kq�Aqa�J�.�09/�fQ:5ƽ�CT
,�]�_�5�R�|��Q�$��:���c��܌|�e��P�g�+��\�w� ^Hh���І�I���ZX��ΙEt�zԺ�}\�
g7X�t�뵴�ˁ�@r"OT'5+"�7s'FF9>���9�PBg֘�\>L��F/�u<�O�T�o�ϊ�8�wB�TK#XP�I|��(A.�;�"�}&[���<N��!�"E\)	qf��A��E{����n[�Pg�����*�#�CZ����K�A�߹kjy���x�d�.��[�`U��bcℑj9��O�o�w�b�rP��f�bT�b)�ٺ�����~v�ѓ~dP�Gc�j�XV�VV��E�� �v�~�Q�jP:���C�x��/��� S����a���g�]��L�n�M����Y�k@�ɐ�u+g<J��-�3 �?A��p��g$�AM;�:���kזR����ȝ�J[��]a��i���
�,�ò�����y�2�E�����������a�jQ#�����H��Y�@}BC(6qI���"�(W��2I8P���&y,��Ȃ�IDGI�`��0e(n��Ks���&����k��C�������}Uv��J���S���T��%�;Uy�,�)���\�g2��Ձ���&J�^sص
9�09
��N�e�Y4����v5��Zn��v���g�4/��qģ�T��x�'29�`\�8V�WE��ަm��_[�����/6c	�Hp�	��v��F<<��3<wF>��V�b��6�Q�c�ߒ��M͹�/�IN��$�ȕ��*�p��E���˄̯#{��o����P�N��Y�T�pI�$�EL#m��z9�W�<-�ӌ<vCO� �j^_����?K��d�]�CE���f1f,<��՜�@�W�3-$?N� rc��d|B���0>Y�)D��h��)�晷�4�kie�GY��y�����@�p �	 ����E[��\�T!0!��#��>�F5m�텝y1�������a3c�`��D��H���zɪ��bV�S����;IT����	"��w��W���2(�dz�O�"'��Z�2�`��9V.��Y���Ǜ�oqT��.�zf� m<��bZq2�.z��'��SB�B�<f�$k��z�.{c �mR_iD#X���\-�	Z�v�����;J���R��\
�<̫����� �W�?�X�JJ�8��[-l�ґ��VS�)[W5��Go��rL<�uJ�J�Y�?����ho�f�1����Vj�$�.o�5CTa�
��d1���7}?
�\��}f#ˉ҆��F���<�������5�-0q3�{ؠí��M�RQ�Fk�ړ��n������L�(u�W}��h�BQ0B�����
x�|y�v���lL�X�͔a�窋$��D��b��6y�6�Y������ig�%^���xNm��. v:0��5&뇹�#�T��Gb�
��%�O��J�ݱ�d�gG��|?�$�b[)H���`���������έ��d^BI�����r��]���ÑL��V��=���jj������(d��x^Dv'$���p(	i�ƚ?(�V���ܤ����61��=ۛ��*I~�૥��h!���/�WL"b��#S���AO� gq�T�r-N�s
I[�Ŋfq��(,��;�0r#��r{�/�:��c��� ���0C��^�~C�]J��:����:~�e�DG�����O/҅����v��T,�S�A� �`�-9m�׵~�z� ̲m{��C���B>�*1�w�al6�eӛ�
+�wUA�����>�Ӡ�W
r #�t�������|8���q���-�k�M�za�\{r%�C��cO��.��NH�>#'7,��px�g����Z��(���s@n+ ��`$�뜃�5~�Y���/��2�x*�5HwEw�K�v/� ���o^��d��_��`�:9��9��g0�.=H0��%�B4z5��/
]�"r:j�P���ܬ�M�Iw<�阯\�
I������$�|����L\}����է��X��٢�)&Fk8��ֽ�g��$�2�G:�Mn|
oR�����ֲs={�d��jp��H,E�#k[��q�ߩ���l����|��)��m�>���V_*E�/v�g]�3#��5s!U�s'��-�Ϻ��	R@�nh���t�¼n8�Y��"�����X���]?��w��>��j�����5���ix\��� ���Zn�he���pF=��G�|�'�jk�Y�Y���)?�͊TA�����c1��'ط-� (�Z�o��9`�a_�jʙ���}�В�����?�@�K ;:�xl�hn��"�?��A#�ԝ#u�3�n|<R��ADVO&�j?�|�
C������
�&V3��@/p6��ͥ*��o���{B��h�L�<� ��������G���8`��!��:+�3�� 'Q.JM[+,Y��7~"�U0?���(���U����,�"E,�|�5��ݤ�T|�����Jg�T
��	��A�#<�ǦW� ��C���6��4��=�?I��l�2����=�mɝ�Ȋ�Mad�66�������$������-7F�r����e��.*?l��G�_���*�����I�;7ԉ�6��l�T]k�k򶢘�欤 ��� j��
Ҫ�}l`�a�O���P��6Y؂���v@tÖ?���"�9B7*!�\Ic%����b��t�د��*�cF�H�v�|�	
�HH*�c��TX����Hm�g���׫��P�%�dw��į)�(T ղD�����6�ڦ^�Q����5�a݇rk�lּW��'��?,��qg����!	<tfLܣg��;���X���Aa�4]��J���t��U�� ���-����$	.��C;�kbWq��"�p�TZ�w�4��2;"7sogW���
�`��T��O��'�D���R��k�(EAF���,V��ST�#�cCR���J�Մ|$q��[묢E�����%��k���）�M����.���jq��ɡ����:-��~�	Q�fH�:��ww����@���L�� ���qt�/@��T�L�f�?�W�GL��v��2�2���l��3�#�_��<*��1f<�9$w)fa/��'m]�U����p̵��C#͆EN�$J�L.2��"+�F�<�6T��	8�|JO!^�m�)��`xf�%Uӷ���H1[��,�����k4�H����8��y)�-�gR���K�ê=#��͡�bo��[��?�C�E�ũ��\�٫qm	��ZGQb�>�5���$_�8���"\:�L�؍�钧2̉�[�Xyy�K�P�k�HV�}`N4���B���6�/%ZA�rB�z4M�����b_�@Gc+J[s]4S�9�퀌��x_́Ҥi���s��%�� 3��5�<���Z>k-́3�|�Bæ�7DP�e���`��I�գ{c>.n���tO��az3��>��wE�V~q�MN� ���!J��4C0�PBF;?�K<b�&<A��0����p[�H��F-Bk�����s�މp�W���H�f����Dȿ#�؆��?�lvi����E=��Y�3���El>�g��" �b܄�+F}�N�
Z{�4kYy�
ܝx��D�d��߸I�t؈��9���xڢ�Rc^�!��͑�M;V��6�sRз��a:�&j�Y��Y}����<K�\Qo��3�-�?�����j��(�9��݀��J241���&l��W�
������Cd������WQ�\ź��w�}�_6�k=1\wTFE�tC�|�Z�UQ��}�g�9�+w���-X�t��\&R�P�t7�5��B��!��	D]_T�`2��7_L�SB�qS������k�oZj��7l����j(b���eĥ^�i�Ű�,�apЋ ��V�y��C~%L���7�B��"�� ����z��<�������5o��NT��#Iy�<S��U�l�J�frwpVo�ʊ� ��K���Eg�]4¾��X�U�{�[
�-S���P�c2�Va�+q�4��9k�g�(��o�KL{��J3�^��Bn�J���Ŵt�(Ռ~�)�a�n�I��W���;A�ƺ�%��N��]d� ���TSy�m
vꭨPL�;x~���5g�f^2~�$�ZtPk�3��f�&�9��C�eDX��f��7le�;ש��ܐ��3�0��e��H���B{EW6�m�@�^]��Qy�_0[�7�Љ�i@4�D���PyA`w�V�/I�1	B})�R]��+R�u-Z�Q�;,fp�ZL��UI���É��Z�}͵=QR��iQƈ1���7c�`s�U�y�N���+�V�S�M������h����j~�zD"jɎ5�i1b��V�қF/�r�Fh��D�7�D���R�򵩁���?�G��n��HT@扯.#~�̥~8ݿ)��7j���lX!ܴ��Y�g�*���_!^Ԝ���'�A�X���U���f(�2&0��߃]�-%��!`3G=���x��%a$]����Th �-uћ;w=qL���`�h����g���w{Bڐپ;��������x�p�xM���c%���&d�p���iH
��ǹ}gn�Pfrԣ���Ȫ�e�if�`��N�~���&�Ryz��0��3�ǋ1D�UQ'k&��z��N-FC�t�{� �� G"i��e��P^�������R�q�ȼV��z�e#��M��"	C�d���w�HoO���dEmQ��Ꝥ�cn9���K�Lt�1+R�g������y�t�*�  �k�h�Hw?톅�c��(8��ձ���?��#F	�y �w���6Q,���7��k��"�Y��&T������|�%�߭�'��O6v��Í���Q� �5C����K�p㗁�Wjn��;0�C��iK[`�&��>���-x&�� �a�N��Q:�=$�b!"@h���JB��W-&�!"�O�� �u�����)y��BS)i3�qR�Z�����)��3/e01L�ǯ<1�mvS
�d,'+� +\]qy�~��J�:����^�Rz�9����&�k�\���ZUL�:4��r{3K�O����B�hVLT��|V�'�Z98"L��{(@��)9�s��)݉�n�w���!'���܊Ă�Εt�* 7��KA?����f�R3)Q��Ew���L�����������Ǟ`�
�^j0�����)۽��� �H�d�֥Z;�M���`�]e���>]�21����	Y'!�3~���������jrr���-��ftP�c���B{����������1����&�ѿ��Qד�){j��ĵ#:����"���o��'/Z�,�1��
?��!�#Քu�J!���ˁRfc�B7�̈́Ƒ!4�����T��k�|�V������������rF�*��j�5�UH| B}(��1��%"�XLN�4rC��PF�'��!�C���1n��D�4�+�t;gpAPv��A�|��k��(;{8M�A�6�I����D+�Q饤�Di�1��E;xQB��>���\?mML ��pi�Te���#�߁N
���h�f�s��<�&T1�:���֭���$ �Zhd1��g�l��.��h)V���D���O�����U(j�s����7�0�:�z:o��������zd���f�RM!M>����M&��:�m������Z���Ҧ�H6N�`��J��R���a���o�)-k�Q����0�po(|�+��g��T+?�D����_w ��'7���߯��<��Bz��> (�WW�{�R�;]�H%5���<2�8�)[} �c���޶��b���飒sS�΋��89��^|���q���� �)��U���B5N�5t`�.mmz-����˖}���U��#�~C� �4�8�T�.p$����SYg�*Ʋ�_�J�����vov����B��3(��<�S"�w�hls������ں���-�)�͑��0Iݤg���/������LBc �d��#U����5��g�%Һ���p ��DN��W��I0�=D�G�p<�_\*��7�@9��+b#);���w��C���P2���t�uO"�Zm�^�8�����E���Y9�;ɴ):�sce=	eq�O��7�e�{�AA�꓀#4�m�a2	w�?��ͷ%�K��e�C�C^���@���ɫ���U���*�H�[��͢U4|���d;-0~�`����H������ۆ�h췶�����׉��\4��ܥ fC�h�ﹽ�P'���S��y�[T>���f�Ӂ>�S\t�}@%���Z�ָwX�f�P�TՋD4�����Bl���2�Mq�p�&�\2�萹 �7(),~�sD9� ���Y��WЊ���)W�/�bn��#�_Rn�~{��@�Ԝ���4�=�î0ԄV�u6�jyy-��af�ȡ�g��_�޸�n��ju>������m&��i���`�kf/S�@��J
#✕�����U�u����?h�t��v�g�0�Mx�e����y϶M���	���B��p���#*!VT��ҁUΔ�pǢ���G�aQ ��֙�/�-��BV`ep�����ܓe'K���[�=�K�%z�t+0�m*'1���2aJo�b������F���D�����=�1��k�c�ϓ#*��zI��5>d��0; =�S���h�P�"-�ހ�u���S�T��_숼$Qt`$�oУm��-�g�<�'Z�a��G�ϊ3��"�S1�=;����h4f��3:xA�wv�t�؞��~�܋lr�CWd\l��gs��~���_��L��ÊƏ��yF/$� �:��!�Ӟ���0� ��,
����I�����V���2:�IZb�����g�s���q%�D+!���z����������)-��w:�8+KqX��Q�=������/��ո��dC�9�`��"��@�����T����g�R��`x���w������`6[��"�������f�~7+�8�I�/�����N�D�x�c�L�����s\ȫp'��;G�gYgs}���p.j����mmM��&D����:A�R�V����'qY[�H6j�q��9%����4���k��(^�W���:�x�/k��!�ڜ�Gy\脣���CI"H���8���S��7�V��d��j���T'� n��7�-� )��?W�|��l����T)U�?;(t&��|�j�Z��4Mg_%�b��8�~c�F�������_C�Z��t�V.{�,���b���rǨ�m�������Ѽͼ��n�,%q�H�M��_ʝ�R����;��y9�Eg��(� h�|{��'<���\(<�?����{j�
~��
���p.]� F�V�Y��S�B[�vJeS���ض!q�bw�w�x�ݍBoC_�r�4�A��B4K��O�d*"��A�ZwѢ/��gp�V⮬R��8��~�8-������
�R�$�qoޠ\�y�7��'��*N��ޑ�[�-�Cj]�Rf_���)��*��M���=9����$�O���Sȼ�C��f�e�Ҫ9�wJ�D�Ȭ����LI��a����@�����^���-oC��:�Bj�/Q�goU��IWɚ����������v>
�����Dy��Fy.�@[�|8��/��S��=
u0���'�f�n���j���]��k���A��t΃M�����A�x��=�g�q��M���
�da���x7k#�,1}����4��۷hݍ�ڇ΄	�j���>8p1Y���)�s����ȵ�z0���W����<1HA�ݻ~5L�/ܭ���}�PYW,�<C,�48�҇9�@Y�j�V$6��W��H�7�t�}��\�z�b�Hg;����2ifB�$��{�y;[�a ��"m��I灟9��x�^`;�>p�����P�weJp�܆�A�D�T���]K�f���V
�0ԥ���F�1�l�)�����]%k�j���g���<������{\!.�x�?6*]��l�r�� �1���1���R���\QHͅh��>��
c�.9�ĠY�q-[`l��I�@2fF?S^��������WD9�m��1���(�����E܃��*CSK̬07��R�:?+��� (p�3�#�J���H�W�!��5��3_�S�&k�ߵ��Yu����[DD$�Wlw�µ���fRZ�"�NljiI3���ܒ��h�H!���k�N*^�l#����:f0�@Pתk�F!$�wY4����q�[��(�H�Q�L�N���̄/��>یj/�Q^gX�E��>�=��ߪ��Xe��}��h������/�oBϐ�Y�0�x3���XL��ٖ�6���%<���l��s�3BhO���*���F$FGX��y*�R���N!a���U�fMƵ��m��k�����
�jY���Oy��x��}p�t}�â�,A/���o��x:	���F�Ԇ��Y��EP5ˠ5MȝJ������9�Lk���HQO�������0ڳ�d�֢�Y����Lx=E�����<��4�q��\��t��zdA�-��s�}�8$�i�*��1��;p=�ޘQu��:+����`���_������e�+�s�%�CB�Uֆ�Ň�	��)��v��N�@��>ᯜP�LϽ����K�JTh8]cѴbθc�V��rI�R�L�'Z-�d*�jb;��y���R����P�I��2��$uGC�绍�R�qz	um����u�l��Oy�$(�O�5m� ����� �k��YIKYOk+��T̣����l[Ce���U��r^Շum<Ĺ��9� ��y*m��5�LQ��w�J��S�K�>�L�_���L{P�3{�'_G흗h������qg�(K�	p�>���8�H�ߡ��J�,��8[��b �#�?�[��	��--�O��c]ܬ��k@��~,��]�ǭJ��^<��Qt��-�	w]��X�f�.9♈�u#�cD���e��v�0ab�r�;�z
�i,�%n�|L�=;xG�<���p����,�"�4��\����v�52C���]�\��5Wb�\�#�c#|Z��R ��_t�y���Ux�KU{�\��ec&�	���K�Ak��r��7�����1��PU���Jp���5�ǔѽ-���x?h|��ૈq�*ͻ���x5�6�(���*;��%7�u��ɐ��{���/�
��9����n�328"(�ſ/�C�v$�VR��Im�cF ��٘���Wضil�,L6Sp���	6M5��邁dݠk����C�����uv�T�s�����hD�{�]{��%��i�ye�2�ś��AFQm̸�#�4�#�2o��s��o}m��RKҢ��k����ŗ�f��r���a\���$a�+4��oC�1�ջ��"��n_b��i�My|��>�/���� ��p?!�%.E)%��Sw�qd�<͐�5(f�Ƴ>��\�d�ѵ�+XB��KGt�)��c��/�rѹ5q�>��\�s	���tl����k��ۅL�HvP!�E��e�0�.����~7/"��]�9/ܱ��ʍe�A~�����E9����@fł������6�s�ar���$�K5Sgd"+��ی�y(8.�q��?G��~�g҈嬖H^v��	;F�qî�[Aބ�'x	8&����w�P�)!Dm�"��T��K�#l< ֢M�\�Qp�|m����C�3�WѪG�o��'J�IY�v�
s�n��4:b��+�l��)��%v3�
�F�(hE����>�(��ג�0ڷ�ɞ���X��|�.J/�=��\�ґ�/�DA��7�'eW��N�2XR�+$�R��ce^��&����R��LV�ؐ�q���C�FDE�5��ޡNgnq���0�҆���!�14���R��7��hϮ�z�
Q����Vr�6������(w�#�sE���M��� �Mp�=ϙ�K�_���� A�bdD5�&��c��`O���e�>�I�J��C�k�^�>ӍҺQg�l->Ԧ���.�� Q0���Kυ4�Kl���>��uk�;�Lk��t���E[g#����X�����f	&�)��q&}z���~!>�d�u�_��p�.����>]ҀM���'����𹆧�:Ė1��x �VM1�%:�������e��<M���i����L\GF[��s�/\�+�3g�.�A|�KwQe��.{G� �������$�9��#�'�D�
��`)����f�闑+2Wg�ߦ��74ھ�hcۡ�P���Ư�D�q0�K��4々�!46��]��^�ŵ��÷��'�/�鷵xw��a=�ii~VK��(�����2��`���Cm YQR���lSx�+���Ǧj�qAL:�hB�RS�����rP�,
��z$֔c���)b�Q�B�_��4�2�2
0�mc�]�ۙZ�/�L�OEoΘS�	Hi|G��tB�������8�.�(
�Zw�D�
Zkia.�v���	�
ب�F}�3�|�#�%�Lf���O9�vԋR+�<*p`3��&�ŭk-��[٢�W2�٥gB���ZOq:W��� �����5��2�/��� �ą��մ�c����;d�����dãh	Ȼ}}-F��o&r��3гȰݽ �'�z�`���I���_�Xƺo�P�_
^-}�J�hn��JI�|y���>*�Ё��l�д���g�Ⱦ4���Y^HN�<Dt5��K��� UB�ZQ���{��Ȏ�?�,_Wk���d40Bڦ�=�E��� �+�b:CjJ��:�YJV1���B����=�*��#r���[![�i�-��&���%�p�V��C�����}��[�.%0�\U�F;�����+�w{p�;ݠ�1�_Qk�G�xH^l���g8U�~�S_�P�@�Ԣ�ҘO�K�Q������Z�5?vp�i�꟏��M�I����u�+�����Y"[7�?G^��^p��G���s/���!�oP��19�dp�k2��Z�L�7gv���"�Vm-kFK+�����ۦ�[�k4!E8�b���uհ=��%�Y�/��֯GbT��M$:	�zd��aԍ�J0�J�.َ=����5�RM�~����Ƞ�z�\���r�>����L�s|�>���7��hg���>�hXq��R�2ET��Q��m�N�xA<�<,)9�5e�
,��p�¸�J��%�	�Rb̟�r7��hE���pF���p���=���̉�8HB�
&r�a\����E�8ՂүG$w�I;���57'-Kq9��ഀN��.xF��|�v�l�����p1�C0o����Y���������R;W��8���Hi7	�8���� �>�˜}+��	b��--y��<��3��#�^��[�C���[?� !O�F�S�&�e���� �B� \_X����y��ѝ�n�А:�+B㔉�%���3�KZ������XZ�>]��I�v1oN8��G�]�3�#]�B_t;�:N����k�0L�X�/�<�:�w�C�DЬ�{Q%�����.�����zA|Α��?gSl��/�{��B����B�+�
Bn��~�?�"f4q�Ō�����F�Ph��gX�~�|����c���f��_]gM���P�;�������3j�=I-<��q# �F��F�[��ٹR�ஓU=��L���G��.�/*��f09�o������q�=�E1	B��=��Lg��#=l��8����t�EI�r�A̿��b�.�
^���
�50��kԣ��~�EYg�	�\�\9��]��qAc4�B]����ݽ�B峔@�3ʜ�$��B�"	)l,�=ӫ��|R�͔�G'�~���G�<�k{���b��P����P�0��'�eU`�yE�3��$Ė}�w�(U�!�p�Њ�kn�E�����U(��12q�aeO� cn�#yù*Dm�k}4����C�Q�jR6t ������0#��&���W��!nm�3�k���S���b*i���^G��xf���B��M�^[r�Oօħ=5�W�&c��ʳFh��������Tă)A��y�g�ƅ��&��L�����6�r"�����
�-�O�82=��;�Ƨ����!���
�"ޕ3��ƴW��؏�:��\�^?�b��q���\w9ď3�êd#�]>��N��P�ߞ������ޘ�O�=�x�t#1eֶ�pr�D>y�ڿ^�����t���,���}*EV����uRiS\ݖ����%$�����!Db��H�qf��	&�}�5�?�ZR8�/�@�k��v[ϼc�"6~�p���O�H�,=Ȟ�S�b�d�1F,�e��C��*�ܳ$з��T�bgٱ�Ipe��1y����V	�Ί� �)*~_V=���PA^u�#,�\�8�)�oG^��W�{�Mn6��l�''���M`��%G&A��iH�A�E���0T|?ݑ�ǣ� �bax&������4+��/E��zE`}�������~ċ�:/�Ѿ�c�B��ڌ*���F�`hY�>�V#ށ�HPV���� $���>��LFAoO�BX�G��6���8o��gs	�C��;��N��	ǃ��h�HQw�=�g��m�6b��Ԯ�@�[��(
u��ޒޤ���ø;�&�8��VGd�d�Nf�F�YixT��B�L�:�w{а�.����b���|�t�oAr�o�Y�_�Z@z��X�ێ\1�(�/��%���9�N�)$���-�]0��Ĕ~��	+���ƚ�����!sӏ��t�>0��U�X4z��lV��|���LcQ2��G]���/�[�7�k��;cl��~Kls
2U��	4|�nJˢ�:L�)bV�f�qv/}��G�JT_Rj+IxI��5��&�n)(��-I�p�e�Z�e�n������Ԗܶ�#�Ү��S��C}��oB. WkQ��A \%�CZX��#����'��r(�f��<p.�;_����m{p�R9�gw�/Amn#��hJ�v(���Tm0�V!�\�.u���*�o���T�P�gz�C��R�ȄH�'��;	�8X��D둧t5��e�k������b�({ʖb*��u|�/a�Dh���,\q�i:r��_�>�{���i���P�xtݰ]>�<��e�%��	"���p��fZ��5�+���[�cxIiVٚ�Ⱥ.�Ep�� �$��0��:��'{>��3ZGs�`v	ώc]�Go��'=~MVg���Л�J^J+Ց@��N�XY&~�z��Y��.2�Q�3/�|ӳ��TeMl��U}���t�^NRfC�4�����W�������[��Q���>�@
����V��(i�!t�r0ET���M���j&|֦�#�9�|K/�.�9����
�@�gZ���-�cYs�L@�UAuw�%��I>�3|s����!��3�+�_�D�h��aF���y��)��Z���1]�Ba�sI�4֔��@A��� ��&>;m6�ȵ���[0_Pn�����z��s��.��z�����G1xK?�+2<6�3�h����Ɏe�#g�:�apL�X��\��zP�&��gՋ�����~"�(�������\�t��zh����M�ed �I�����z�L$��Bd3�Aq4:����`�.Tդ�W�f�M�U��B��	�!|��y},��0	�\'��òP&&��RK]�жB�a�:��mDLM�{�6�k5�k��U�j��B�A#�F�WѢR,�EW�'m�0����ő/?�M�$ư]	��Y4�^�g���r{��;��֚�D�-���#R��k���M�t�!ʺ�;R��v�8�^�M%*�+�I�1dp�"��+��*9\0��4���c����8sT� O۞�/k)X���T&���[�5M@����w�cD��@R>���]���0M��k�<M����>�uV�v݈-��N�Z�M��AщfC�ѪHδ�?��X�
&��a��e��$��o��oQ��It����ޓ�kG6\i>S���i� �wvTA�}�e�7l�a�\�`�\J�L����q��7��ݵu��҆�ï����g��C"[i��~(#,�b@H���B��_w�Մ�tI"Ǘ�ܡ�=��N���J�l$*"�J_�N2�Ea:�o�A�[UWa��(S��"!�3m�.��:����N*tΦ��j(�ڝy���;<8���W����?�򵧟,����3�	2�=_O�3j1�٭�����F��0���kd�޷a:�6ш8���T�(<���7C\
��|h	�Ad��A�3��
�P��2�t14ee2�Xt�����S���(_�7�6�F�j��ˊ#�|��`v��Qҥ� 9Q'&
���~,�D����ՅGG�Z��G\4~�����Yb�F|�2���7�a]��x멕,g�����.�q� д���� ��_�%$��������z/4~��R���-n���o)��x����x
b>�:�.�M��rD���X_~D��B`�|�L*��X�<�U�f0J���|8Ul�l���l�ðnl<�Ó7$!�e��{�`�-���^b�!"2s�@�c*�٣������m������3hBL@����ņ��⑚`��Њ���*�˧���!�b��s� f��bv��aw�$i ���!�<�ۊ�s�Tli�����^'�흚�r_�z��9k�`a2E��m�+� ���P��"=���,km�r�g~R���d� ۄd.��(k���5�_}��c+1N��R/^�TT� P\��3�Ӊ��gV,h�6\�4ԶE�ɥ�C� �Hd 	@U������Yd[^��"{�CYH���$�Yx깚���Q��B��$�� w�\�8�E���=��d$�A�5�Z:���� M�Jޙ�g�QmH��C��0����nj?Q��o�;���\�t{pҷ��bz�]mҮ���"j��>ҤӶ���Q;��`�������ߋ_ 8�:��S�D�ךC�K����<AGPJő��[�8���A�Bd�bޞB�tgw�n]/�ܿ��F�H�����\����J��/�e4��#f<֯�e��RS�����y�=��R�yĚ
���@%�œ�`���Y��BA���;�M�}�жj#Ӎ~q�7�Q�^�AM�c\g֥&f(l��);�`i�H�)�e��qa��o�]]�ɔP^�dm3\�#4o�}�KfF����{T�K������h茅˃�s.�l���� ���<���#�4Q�"����Z8�L`�Wҳ��IX��!��C���>R����)�a�����']$�W���4W��5�\{��ҷ�ԸH�T�F}o���H�$��55}����m�7�꜍��H_����4����R��<��*��(e"�����əlJ���Ϋˊ}������tRvV2�<���:-r��<H~m�~C ��tH��!g���_]�b%�T=�D_c�c��A�cM��ݶ!�=o�u=�]ʠ�||�%�o:C��=�|� g)��6�������G�L!�|�]�����xҵ��c��K�
vlW,WJY���}u0A�+o�J�~8bV�@#��I�G#끸�.�S��BFO�FYuy�<���TA�H)>}''Y��������BӖ��^��6�~6C:�R������&���r3dS�Ҟ�������]��o�s�r!�঵�^�8���з�P�R���M6st��۪p�2�S����,-Ӂ` ݂�c4���ب�	2m�c��O��l�j�a^�_mt˩"n`1�G��e��o a28͡�����0���z�+�\O_Pm5):�G�=�z�Y�ćC0춯�7#P�\kg���K�d��Jn��nd�;�@'��̡u��3@�X��td���S�0��N��?��_��
�>�.fp�~�X����JozH��씚����,�x�O���hd'����?T
���������{�/�~�T�D�3nl0{,H�{�_�"�#3�����h`m��F��4�? a�>�b��\�����j��n�i����5p���B��G��0��)�O����M������O=7�&�F.�,e(2atڱ������A��_ǥ���v�WU)SK���GMm�R�����Ɠ�c` k^tw��,oҹ�$�x1!Q�u���+m�7�3l�*���r��0I�h_�)��@�@�	˝Jo�Đ��������i���w6�M�Nra�4��`�i��eU�@�:�+�"�{�TI�L����ތ�F���j,�wv���I��6���={��lEE����bv�k�(h�pF�~��Έfft�����l����P����Q���p�2��	+���})�3Sg�W�&T�5�W����S���&8��_ڊ("NՃM��L���M�&()ol�<�O�+�v��t���b�%¸9�R�1�LG��U��~w������(y�P��u���{SW�:)zk6�[��Ұ&՜a��M���m��1qA�ss>�lE�zF�
3Q�ջ�1_���U���>]D��`lZf�A��}L�	�D�	�jN�t�Ǣzg�I���ݕ��.���7���򈔗
�	E�{�p�AWC�ٕ��<�-���� }^o���4n�8���	��2��Ejjm3����:sŦe���X���k�l��d��ؓHU���j�����C~:�D5��U[��� �|EE��R�r�h)uŷ��B8r�	��h�[��o���F��G���>�rL��h�1��C4� ��8�r�bh��Ӝ�Y����<�F�GHۚ,���|�/8���芽�n7O�"e�Ia����ͻ���^h�Z���.&���"egKO:z"k8�_�t3����f��̂f���K��C��N��TH-�q{ƥɼb�]����o��6�#f���!�{��t*[�n��p�������j���.�l�4�~��bR|%��J��V;�O(��4!�9�m')��4hr!Y�I\��rl9�R3���kp2�-�ӣ84_{��׀H&���K�/e?��0�B���ee�ë���x� �`1y��uD�S�e��m	��OmF}��@WE�mMY܆,+w^I�d�l�1=��M~;*fP��|� ���~C�	�sv ���=�~���"�ƕ��#�g��eG�Z���N+��j8jl�N�6��0�I<�VY���0:M�ꙛ0���D�c2T �نz�_�K?Bv�� T5�&��8��6�ʂ-�R3|�8ڳ�����D�����}�t��ݑ�,�������mP�)f/�L٫�MXY<�@�(�R7��A{Ǥ~�Nk��N7����ͻ���a��.���'���N�h�IZ��s���������Y����qs�������$����6{!���T�3��+��D%�E䖬�nߝ:�ՙ���:W,܂۟i�!�)U�n�'�`�;d���V����_m��׎����������/~*��*Y��0��6��x��'�H��CF�`�q�����ˎfgG��G����[R52<n[�,�9�����l��]�g��@B*�+�4kr$��X.��r��aq�QhLˈ$Œx>�f�4� �����#�'yhr�O���=�c�A�>���(b^��x}	_eyqe�	�p�#�ጋ��SG�tk��5C�L�w��	�^�`5���zx�j7
z3���J~W�ZCJ<��`m�c�Y�A�P�[H���B��}}װ1���,cqɰ��m!��?!8��T���+���q�;��*�a8ʾ7D��~JS�mp^�'�Wr��
�	�m���Wf�/`���N���"�T\���.�fo��V�9�6�Q=%�=��A���J�RJ#�I��ϲ�?��a��9�^�������|3a��+�6g[Fre*�;��Y=������0�᪠*"4A:�y2L��l�n�5��Q -2��Cg��� h�Kk����!;��t2��W\�Y���o��;y��R�YN��ܪ�XP���,'�S>r�;�c5�6��'�٢�8䵍����t��;����T���Q�ra��+���-
��4A<\�f�vܐBy�Q`c_d3�X!c		�#�,�e�*U�G�s����J$����t��r���ϫ6l&2E���/ol4<-���V�lz]D�r#��C�3|��su�^��P �$%2�iK<|���-�m3�W���jX�w�c:_*7�]¦}�S��wJB�4q�{b3{ז��*��z9�Y���ة��`V%���T,T����'f�k7��@|aM��$i�L�g!%�쭃��Z�e�n~o%�@�I�B �"�>%���7-1��2J�q��Ηc������ň�Y[���f�a%�Z��f�0ٺ�����'���Y�"l	z3�&!J���9�*ϋ�{����&L��0Y~Cr��T^-	-���պ��&�uK,�~������5�E�cɥ���u����7A�]L|�ӻ��),�6�
�:��-WIT�p�|�*-���u����4�x`'�"7��Ôs�㶝�B[B:��~��=�=�������ӿjf%'���Bd,p:�� �hg�����D���T�I�MW����{eQCY^栠��N���� �0����vz)K:B�l�^WqJ���ZH=�{4�s.Zn�4m�j�V�?^g=׻17\<���vQ*��&V�1�hs�����WyF/MǙ�Z�4\�.L�:�ڄNo�r�_���%�~:��6]��TQt�SFz�CE{�c�gȴM9[��S�B�+��Y��B��U���Z���u_����OBBq�un���ع��D�'2�̹�y�R���!W�ɞ�c��nL��<�##�5%p�����s��E�J�� j�Wm������T'Re������)Y����<��L7�(��;d�s?8�pš��!�����e��y	�u��R�7=���("�:��n� ��k�n�
�{0���z6�x��D��ƛ��w�e�T�9�e��S��}�0y7Fl�����'�@�A�ޱ��(Y�8��5]����óQ�$w335��E%n?�_1C�����r���bK��h�-\K�zQ�/�1���ѤN�͕"�6Q�U���L�=bG��E�[��f�V�/u`^�#6l_��P�q�T# 6����OL�����9
N$���̅K����β腓��,����70�h��l���ZY���q�`fm���$ߏ���A��Q���Wf�/喟�ږ�ɜ=��[����z2G|K��)L���HH�b]F�ш;�|�pqCWL�)�L=�i(�QC�h�1B��@K������ycw���z��"���]��xٰ���u�s �Ŵ���a"��2E�H�b��w�\�1��l���S�����qf���_	�6F0c�f� ����������5���� �dh�E�t�R"<,و_
��L���`����2�̊ȏ��o�8J���a�hZN?��U���l�8_נ.�[���*�8�&;�u�8F��3
��]��x>�-�f08t�P�?4&]R�a���[?�.�Z$���9���Cy��P�I�;���"����	�J�s�ɤ��t�b�Jfppw���QR�R���I����+%~R�<A]���@�§m�����0�	���0H�����"�9��e����O=M  a� Tј�u0�eu��Т�B����k9~�H8���;9�pa-�ҁ/[��U���٦w:Y�q�jlɣA+_B��[�Q:�w�~V�/�fK(E���O����U�9v��%���X�ʎ����n�.�L��2� ��,��=M���)�mP�c�/?W�J��>6"��NP�����Q�*�fX� �Rz����<oq��sNm �'?���V��a�C#4��1����/����Ӕe�Q�����:�.p��G��3��/׵����27�Bl�,�D���M�QX�0��Bc�^<��m4��35:@��|��4��kxA�0%4T}��%�XN��ѓIY%�m��᷋,J{����޽Qew}�.�go���(�=��q@�I�ްE�#�~�-�x�.�:����dҠ�y��B06�R��/�B����	ʇ#J���ix�y�y-�ζ�鸓�}�
,�B�5��TF�a�;�5��+w���f�7�k�f���iX_��N`����"��+�M!���et�4M����g znU��xȦ�+z�r��=?�Ճ᡻H�r�ƀ�΄$�3���� ������e!���a�1�L�IB��b�@A�8R��xQ�K�yy���?-g��)��U8���LT���k!��)���<��>�S��<�e�.4�j������6�|� �;E���z&����$m���+��n5�K�D�#�����ŭhO�̼��Hr�.����i]R��`9&C����3��ȁ�����֯ߥ^�r�
����C}�0)/7�x�<�2込�?��o "��%lBj��6U��S:n� u����,Cc�ڭ�Z����3t��}��j�]y����2F.�٣��|l����-���dW�m/�p�,�'����CLSz�=zjKR#_��x���Ѐ�g�:�$�֬���o8��~�>�Y��U�%�*&T�,�>�Y�7�r��O�F�j��fF&��� �c+�&l'�s��� �	��N$x
� qq|0��q*l��8f��.�Y�+�rh?�\�D|����랒\��&we����S��4-1�c�u7@Zo�c<g��-��KT�������x3�\
�p7~�P�P�]i���L�R�=��Q��xܖwC�vZJ���� [Q�k�|I
��V�ǚ�O@�h�/ 	�=�u�d����巋��W����i.�^�"�����ci��g��l�z�c@Z}��VH��ǳ���E\Rh����<&�����j�?���
V��)���((�1�� �:��7�׵N?!G����]���h�].�w���UhS�m�鉀d(v��V
f��ˇ2��G����U�v�1�_V ��n�9�����W�BS� p����b0ѯ�������\�b��߄�Pͽ�r��uܻ��|�p���	`��reQ�i4[�F
��̶TW���j�jn��(�5Q�'}���-�M�]\���Ój����m��QNU;-���Z�Zf2<�g�1Y�(8��9�JyՐ��tqR�7ۯ���,�K!��(d���*�T��W�����G\*����Z�0ѻ��P��po���7��=�f�M�q�%䐞q��ދ#���ң�jy�
d-E1�E9��q�l�()�BVw�+G#!�z�Ѿ"��-��Y4�3�9i)]3Ϩ	S��̩�g�|=��� >�'}����f����Y�Q[Aq��� r��׵"��Ő�I���]����ˇ�B~=��s�XHO�G����U�%���	��>{�7A��[�|�\�>&~0o;����jQ��El���<Nē�F�BN��K2�zl>o�?�A��g�Of}]���X\�oA�����Դp �-e����ͨQ�V��+��÷MI^hȾ���S	&�?^ĭV�b��e`�p���g��>Z����T}���3Ϥ��'\��9�����;��_�{���es�
��D^'Ǽ�r�������P��0�Wؙ�'mb���c@�q����BWh�0��9�|�}��B�H2�`s``u�J���X���j���f��}S�f:>�(����j�I�U74�$���zA˲(�D�B�h�%f��-�9��Zpҏ�����E�0O�Ѳ����Q�́v)�bjW�.���%�=<���{:�MLqG�y��(1�H���1���n���I*���o�~�zʧ��\A��9�G^$D�}��1�ClI\S��5�Ɩ�0^���Y-p�l1>ꞿ`6�A�a5�����h 6�{�sԢ(B���PI�K��3�S��&��[�< ^ґN/`�k�t�����:_.��uD�2D<F�b�4����75��n-_6�����TsC����GH2�F�y�{-��TqP�����!�)`al��� ��Sae�˗j����I��������� ���/���J��5�q �b��*�}(�̲/��ʧ��'=�K���d�>�BaG �I༇��ЌG�I��ٔ|��E��'L2t�S��z���p!��[iR��}}r����AR����Nj!�dAp�_���0��:TT��Y��*�>(���)D`�dQ�^���m�|����+������mU yw�
F�i)�;�6��&�v|�p^�ǲ?J������@�NR2G��ۇ1�CibA8�!���kzcx=q��e?�~�O���� �N�	}7(O��н��v�B�cw��
��?U�+_�T0+Kh�Gbx,�tf^��֡�Î��1�iF�D,�X�3gf]�~��G
�պP�  E�gDms��ﳜ}�!w�K��yҗ'�]~?_^yo<�⿕�&7Mb��@1��\��+�.��X���y�$Eۘ���d7�ކT��	v(ˠ�#� �z_��h��v�)���2H�bY��`X�E�)ӈ+2����?n����
���hd|�Ӹ��cw�e��z�g�4LXO"��+�Z+�l��N� V>d�R�j�fka�ÔOu^����uL8��kL7���:g/�j�Ҥ�	�G�1"��ȁ�"��o(=+��^�@�z"�.�28K��+�BbaW����4��Yu���ڴl^ٍ�;NM����~���*�RZ��]wJ�}�b���W�� KD�u:�َ��B��NV8�Q�3M�9��>�{�G�D�Q�ܮ
6i	ݭ��@yߑ��	����.
� iF��2&?u�9M�4U_��;F��$�i F�z����k��v2�t�S�K���GX��痒@�X6���b�RkƁ~Ybo��${����Mw'	�sT��A��	f��l�m}���nS�pUQi�͉f�U��f�MJ�*��w+kF]�-�,��;��ec-t�W ���k ٓ ��D���sRW8҇�H=d�}J�ݰtU�S��R�	p�4�l�*9">�A����X�����%���MZx��L־�Kr|ZrI߷���6�=�Nv뮈ʻ3ZˎOnk������.��2������u��cH5�/[�k@�ǣ�����<���>X$�Q��{>-s��A̎�`�k�,��!�q����H�m�4q�,���#ؗc)��H���� �1��:����$��G�s���by��382@.�6ե�`��tV�k,;a���i���f'���OǛ��(�Wl�F�sR]���~�u�<�nJ;#$����� X��9�޲�	Tl��G% '2��Θȿ���EgV�5x�����;��$ "��0u�q�)O(��l�������
��ࢫ�a��闓��
�	/�mW8M�0j,"��?廞�鹨��
<��̮Q-I$���t++��W�U���1@��҂�B��G�ڵ* [.�ky5��fzT��`'ϐ5S���>q�*�o,+�;�Ӽ"&���e0W�W� �Q�;)��"�srl�����!��R_>14�����-jg�i>C� |+=qdd��6��K�`T�ʄ2f�B��dED�*� �٧��=�����1��'�r$�hq��q���W1�m�ھT^[�T
]<����N���	1�^�Kmj4'�e��3Tr�ܞ����g����V�և$��z
�m����u�+>w�9D1G+��as]�t�����Ї'xe8��lvP
>��2�ԙ���0�riqZ_���71�OĮMhqs@?�QF��ϸ8@\��A��aCB�����kW�q�+N8��Q�+B?�(;"��ǋ�(x�	��z~����4�A��qɰ��8��nNQ�^B/��o�l�>@�P+d����lS��b,�M�����r�7K��z3XkB��إ�.[8x�k�����Մ2�N�1��j(�aj&��=��";&��G�!�^�q�q�ъ�$A#y��KK��5��ػ�{��~�n�U��Â&�^�6g��<j����aqZ�v?&�gF�i��#�m�K[� ����kh7�Nv�,�����{�"��W���.N�>�)˃kn�\��7���X)������CI���&"�}��
eU��9���gZ��f�����&����M�P��f��r���Z�]F�fLm?\'�Ѹ�\.�&���uWT��ϏDi� }��s`յS�(����!uY(�p��f �#�o��,�v�p��?����g9��5؆�t}��lỻ��/��}=�`09e4����t=����hM񗲕��?��9�+f#���mL^<�{?.��~�^��P���t�R�:�~�sH��~B���x���M��/�ʧ�c�2����r�fL-�VY�xSeEf��������2*NiF��5d�t\��v�Ԑm��^��S*kb�Tr(�ݹ�<��K��3|e�o��1-�8f�J�&�NMy�V���Bpz����h��ȥ$�m�;&E$����j����p��%��-XN�b�^8���,�.�MI^�s�\]+y:u�Z�O�#��O,KГ@m@N6��/�+A����� ��ʔ�f���!5�ӣ�՞>�����]���#�T��i�o©����{[����6���T��b W˨���ʍ�Rϼ��E�#&8V �����lf�&��Y�ēp?9h��8X���ѵ�q���rG���B?HQ�:�ibf��l�S��꫈�uG�$�9ύ���M��R�܊y�w����b�]����oc7H�A]�G��Ԫ�Cp�Or�8'�"��ŀ�
I��?��a�kBM3��f�TH/��UuxT�/��aj�5�	VF�܅yQ��־��H��Z>KOT� h<��^�v�u���PY��4|D+Fڝ܋mo���@��V%�K����: [�M�,�?�2O��x
��8��9�%x	���Κ�.���>Sgu �(5�K ����c|S=:�Qh����ty�C������U�q�A����_8Ԭ߯_�[�o�}�(�v�/�ۨ[|}���,�S
���Ûf5Y9�B�\P]]�$��L�]*0�Ӭ4������E��_n��D����� �j��Eʀ��w�Up�L{�E��2��t��Y&��ǿ�
�`+r^�m�/��z%�k��U)�%��&I��j7����(����6����:u�#;9���·���0��ش�d�y�^�IT�䇙�3 e�s�NiĲ�1w�(\��nu�����k!�4A�XO��腒���`[�)�h#�t���x|J�ō��������c�O�/�M�d�<a|�߾��&��3�*��z��z�Yc�K��6��ܼ���˝,���^T����f���H����>;���Z���mB��3���+����P\��j�6��W�I��a�D��v5�eϋ�jR�T�Ot'K3�gR}���W���R|d,=/��ҫ{��*��qn��SR��<��x��f}�7�y
��J!�Y�qV�ޱ1����=�7�X��S|�	��f�$*tQ�����1�_�c1���֣D�F�1KH+;�I��T�e v��)��M������nxRH=���#4/���dD��Ms��]1?I?J�6�� c�I|>�f{<���	��1~�L�$I���PWR>�k6A)Y��T\3�C��b>S�J5��`��q�#M��*�d�@qш�-��!xə+N+�{=��^(BX��@�8�F����q���1s�R�=�1*r��1bP܋LQJ޹��4�ȞNҵ;qw4��`	��*�Clۣ3�e:+�x <�ĺr��Y˝�����iɢ��� �Q�,3��phU�P$�|%����{�$N�-��(��S�욹49�dp�s��;U�n@A.��zDf��7�G(d9o�l�Q,'�W#���M�F��4�4���V60�Qb.n�5�i�LɸEJ�A��/���QX.���r��J�����a3�FI�K3'D�,��LyB���Y�j����z�E���ق8��	�Mm^@7ߩQ���M�;�m����	P^�9@֬�ٹ�F���w�A\$�A�1����lh��n����$���a m��?�*f��2��1��.��3\�.��0�}���Z�/5c�)�M��jtM��*.���1���M����ne�� :!���y�oiSu͏!��hUz *�x�ȩJ�ѫ�=�i5�(����fW�0h	1!MŔ�weȟ�m�sK��k��۶߱����hU���ֳ��,��w�/x4��!�����'ǹ���ٕ��3M�=�V�8�SX9,�n�����Z���8�'�*����ZMEd��`^H8�~0��0F���@,��;?j���ct<�H�No�t̮�Ѷ����\���KY�H�!51$�a�܍_0�D�5Kd�,�u�R:��I�ݕz��^P�2_���G�V(܍T�8E���`/D��)l�{5Њ+��Іȩ���Z�Й|�;��=� N�6�ŚL�y��6�A܏x(t�$i&&#j� I�u�2��R)2��oDk�4��u��e@.�.���ϐ�FXț��)X(�WY��w0���;�G�TX~�>�eD+v� �w?<p����>��tR�6q�Ez;7d���ŗ&�Q;ʯe���5y��V���fD{��6fB���l��/150����mF8K���\~�%��~�����Z�cQ�����<��:	O]�a"\�2?���m�U5�#X��o^�֒���m���34��|��3i�X���p�$�%�vCr��|���(UK��>+��H�%vz��q�`�]7?����z0S(AV��t���5�-��qaS?�&D���1����	�y,_WRei���������n�J�#C�����(y���ܹ܎��j��K1׳�\/Q"��g^��0��ҮR޳8�>���A-D{b��fp�t�����7T:����+�h�5�+�am�7�0�x_�l�e1����EoE�kJ�{'s��I��|�z�,�]?��u�}��1̦���9(L�P���+ۯw�b":
ѫVbO�x�`��ڑ��c���%�t+{;
��4}	Hq9�Y�a^��'롉���@�8�m�2�[�7|��/M�X��Cd>Қ5� (�9��T�r �u��	��3��H2��p��T��5���mq��ʏ}g���kUa�M�ր[��6ڄ]�����X���P���-Έ��؟vi�-x��[1]?��o�?��e�Ɂ���Q��L�S�g���/�
��h�+֘��j�jӐ0#ͩ��P�lR���BǮ����sf�C��o�< �Pr)��F;���g��8��Č���8���k�U�$���,uMA!���(�iHu��͊���h�"}=�1��N�O"�ѱI�V[�!�!��l$+�駨æw��U�T�}��}�K��e��f+b�"��G�ORi~1��R�B_�?W�O@���:(�O��@���^L������C��Yd<0\��dFP�4lD��3诧%��=����{���Y\������1��Ě~�ĸ����Ǚ\�Y1N �A��![���L����Ug��^���æ9!�\���1O��}[�k����i�0�<�����Kj�{m����7������ɚp�O�VΊ���Nv�	z�(R�S��tjr��GyVT��y ��:�d�zM�G�	H��&؉{�Jō�[yV<�c9�����o��&�H)"N�g����`����lm�7�߉Dd"Y�X��`Tkԉ3�t���D'�m���/��C吨��?�ub{�.ڶzJ� ʋ͝[�$�S��Ყs&H-�l�o��]G��;N��$pO�ڵ�����X�����d'Dةd��P�W��'l��N�[i_ ���&yd�La���LmP��nW5H�4�
a|C���J��=Z�.s��f�h<[5��Ow�F��v��//����O�k�i 1�� k;{��G���55�R�O5�%�	�T2�r@�&X���)��Lİ���; �3��~�QDBT��D�� �cO/�r��|'}�J��"j�
�B7�U�H_����x�f��k!���4$M�b���4q��4��Q�FQ���lP�0����������q~�Ġ69����[v#ج�:BPz�F!��;��s�;<5�Q�1旿x�E{����%_xu��V~��Ӽ�����^��*���/.~�V�(Ǉѥ�8@��1�?�7逅t��er�)�6X�pB"��"=�׻��;����b&�`�*�u��`����r�R����e�<�`L�7K��Q4�o<��q�W��l��D�� �I/�5���&]���&M�G�2{6G�R�ɿ2
*{H�U��n�oc0����]v:V�hP��971�7˹O�Zb g���q����T��N��/9�A3��r�Ķqˮr���sJ`�E
�1��c!2_ۄ"F��!}Ҽ�X�	�����e�D�(�eE�b`Lͬe}Sj�J�
�Ѣ=+UM��fd�Q��	��{��o�^��
����H���؆0����2Y���#�ჩ0�G��"�9GJsWq�@��Y���������<�ϾFc@��*"�R.v)}�h�}0|�
����y�K�p�}��~1��JPL���R<	��������޲�v�KE�Va���9�]��f��d��:Xz�B��)��耂%C������[�ak�j����X��n6E̓ �7���N�&�3u��jL�r���\nJ�6P�%^d�Ki�ح_A��^��&Q�����vқ%2�Q�!��D�G���M�q�������Q+U[I���P���X�zJ�Ȕ����UVÀ
�Wz�2�v���� C�I���U�6�>���.�ؚ}|7(ү���&��i��:�oa��tm�xA&DԵ�B�J`���w�=��ZQ��k��\ ��h2�f��=3��<�wT�gO��r��vqo"t�]D���]��Ɯ5S��5:{[�����l��EAdS���U��fLv��P��E���Jh~�I�"�"�:�X�9@@�e��L(j) �9X6k������cf5������ֲ��bi�d"�8>=�ɧQo)O�[��؍q�;"<X\
Iȿ���R;�&�_US8�#�ySu�����Y�Ic�U�����pj1$z+'!n���YnbC4I�D}į����N�Q�s��!��̭��ǨF.gP�R [���	tE\��|�a�C\~;=�"����-����>ؐ�y���+���|���"�p˙4��u�o.���ۼe�#c�&�Hm�a��>#q����O+�@rL���L%����T�nq��<��ܖ!Oe$<��tq�y�X���'JZ��I���7�+b��?��dy%�/����Q�j�"A��2$l�_�R!@2߿������ePC��̃- ^s�O���!6�@��$(,�<����w�)&��:�����Fg����sJ�BUGѳz�x��κe��)��Rw��k;�I�^��ܥ~�=]}��ʙ�M�9~��-LQ�_|>�)}��%F��ncmV�Ų�-z���<�	O�Z����|�(H����^Xc�{��8��]���^��%�Ђ�В�l덙V|�Y�F�6ي�E�Xf��fC���J!a�rm�)�<NC��|�R����� �G�i��n��ţE���?���g~e�hmZ7��30���U�w�I�R���
φaF�t��?���G�s���1+�W5�7��N��`�5
LSX���@t�l�8���DM�SI�n�����<�X��y��<���I.����!�|b~����i��*���F��O�7t��W�O��*�����l�a��'���V��b鹳$�-������i�#J3���4:8�\%xO���`�h�.��"l)D3�7 ��s�_�:��XZ�{"Z��^����mr�G��6��z��s�Zl�C<�j���78d�R�24A��H�5l�8�r�:��H��70U����1��������#:�=�W7h%d's׫�CVTA�g���M
�M�� ����:�Sl����LQD�gt���tB�YX�s
��S���@ވ��(��.Q��<VvO�d � ]wV����ʻ��ms��=�u�ks0B��$�ޒe���l�!���.�����(�-^m1��\| �2i&5i�����'�=��4�6Dt��Q��K_Q����R�$���<T�{,.Ёe�n�'�6�P;��}�pt��"{VK�k���,sl�сw��(p��k���E�y����+1!sSO0��&ou`/��SD�����}#&̠V�tz�D���_M�F[sU~Dk�I�3�K܁ߡ,2m,���p���`��� ޅ�h�9�����)7�����j���&�wfx@B\�6����W�W����G=����g��4��Ӏ�	&%[(��b�oQ�d?W%@ͱ�Λ5��姰�T���Q�{��)��1v�"�d�e"҇�|O��<W�T��̲�۰b���8��Η����;���N��n�`v�7ͷ>��_ J�\��d4�GI�u1M][R��#tKV��%-�lr�<��L �"$��d����kv�6sH�O���Y�N��񚑺�=�� ��?,kȌ�ۛ�+1f,=����#�-�W�I�Y$��nL�4H��ux���0�@�J.m��)� ޢ��wU��	`���{F�FaV\�\﫵:ٸZ6��ѯv��T#hWeu=h0��7���/��jcv�DnԸ$�"�S�۶j	5�a5q�nu=�y�	�-JL���$`�z�x�S�y0_��o�gL����ט�Q�eڠC����u�<Ӷn���%�R�D��a�aw������v8+����fU�a�Q��M�Уo������DG鿆!�u���K'F��[�ތV	jd�sx��M=z���}k���q���i߆��5e�g��\����Cf��K^_"�����o�2��W����a{�z�#kN�G��-�8�0f!�]����F�;� `���{ƞe�[��tn�\��v̘�o+nٷ��@y�0=�|u�k> �{�H�B)?a]���5�Y����_�1�`Ѳ/��Ｌ�Iq������߫� ꤷ�Y� ���ޜ��o���D9�1�AS���'��+Ⱝ\�0�����O=��c��ۏp?�j�q5\M7�zt.���g�,�دe�<3%��؍7��ڕb)��ظ�sƯ�n!�aJ�b�!���\�^yh�17�V'#�}#���˰��Z�RY�C ��z�D�RAJ��R�A�}+�vgY���d4�����?�SJ�ǚ�5�V�8~�U��O���:��)�a�Ⱦ��fF�x�>���_@ ��dֹ�d'��i��?�F����,o �i"�]��GsQf�����b�т,.M�3�Y���E�X ��[�e��:���=�M��&�ޱ�v��"�)Q�ɭc���Ͷ��|�10�w�[���\k=�вe���ӵ̀ބ�
îTV���+m>\��H̲���9�r��cm�M��Z-�4��>͇�[�!$�s�.��cXP�1�A�@uy�Z�07��F7�gT|�0�
(���@�,N�{�Ov4�9�	�׻~�>NI��)yq&U�J�%�rs��U�x�a�q������U�^(o�������WQ��M��}e�G!�Z�X�>����wF�)[yj���?\��"��&ϡع��tl%�c	��mBd���%Rx�M�� kE[ek�p����V�R�]H�������݁�<�h�I_����!��L�'0�ʈ�wU������<٘3ڞB�s�O�)�q�Ex�f�����H�-��� �r�0�TZ�x�L�l�>}|������d��?*5���@k��Y��ݤL$Òt�����З�î~C���"��_�{K���/'�{�< �����#?ϷPʐ
�m|r����n୕�C�-�#i2w�V��'ll��� u���2u�1g-X����_
���*��AH9��a����*�g�Ȣ���.����k��좌�v�߳�Q=���Q����Z���T��,��5Ɉr_��m|�)��#*ȍ�^��9n�	8��F�P�7zB����
�����fO<� �fY��
�6z_��5��tRk|~���g��SK��^p��2ڗ\G��]�����J�y�������'�x1��h�m�5���M���n� ���@����T�;��Dv�C����6F���2XS������d�f�`
�#%W�,+~�j��fG��X�%��n�@%p\�n �����hC���}�N���T�>C��кb��o�}�eѦ&�Uź5���,6�?�����e���������)ڜ3;ՉQ��:������)\O�ԟ�^{�G��+}�&�kn�<v�xX0к\�{�E�w�5��F��x��`n+j��?HX�!��(�#u�t:���D��~*�wRc��-:!���:p�Ġ$~53i��[���㝵]�p�=��*C������AE%w��⻴��
�a�р��e'��H㳎�P��~�(,�?;ݩ%]��o2.��:/xQ��Y��F����p�HM��G<W�0+f���޴�LVnd?�ۃE܋� Dm��x�ҟf���[�ȡBP#������蜐K���`���zc��2�n���������嶷��qm9�]P�y�+T�.hvO��d�X2��6����b`�=Sa}��w]�S��>�����Pb�B�?����m��b#J���fv���1�fWʦ[YWmB����0��ו*Mx���'��B�"���DN0�N�Vz
LƇ�����J�fiE}�F�T�2O#8��fO�(����
^�s.��+��sA�FG��@b���@�� ���Z����Z�V*����җʲ�VQ(��y��K�pԎ��>r�ޖ95�=����E �^����$K��*&��r�R���Z�j���2o��p��H��H P���*��9�N.q��/ԗ
�cn@��I�׉�������g�;H�f��˷�C"�2���6���4��8o����I�8�Cȁ�:�Y3���8���ԕڨ[��-v��I����dB~����%o(�Bqwlcr1�
[q񢿢����^���9<Bei,�Sz���J~��Z�qq�P�7����Rw�2�Ǚ�naYP6ȓz����HG���Њx�$�s7+3�Æ#7��(:���9�䪝R�.T	e����Ns�,�(����߆�Y�eq�n���Q���'ۻ񠖓�.GKK���z�p.��2��Oj�BƓj�
Su5�l�!�a���z�����x���/����7����&�@ykt����	�u�4-=T�gh�2aǤ��U�K��5+a�� 5l�T�[	Q��"�X[�3U�S���V�b/�a�51��E�r���⺯���n������Zd��ۨ3:�̬Bǂƞ� �Le���ߜ�c�,�h{a��U��E;	ީ9�+$�z`��7�H ��T�"4m��q*5�Yo�:3���"c������A�0(9ǔ��	��8��9���G�
�^q��|R����5͆����L��;I����ɱ��610���'�K��e,&q��q��:�Kw����z�(��u4��9�J�ѵ���<#؀��{��h�p<�l$�~����1ԣ��4�9��0>n_p�zz�oqU^�<k]��1㠝��8���/8s)�Ѫ8N��_�F�6R��!��a{Q8Ih�i�� ��i؃
��e64NS�Ŵ����9���8	�[�aҔB�f�G�g�8�h��"�Z�*����.��]������x@���S�����W]�D���`��Q�g�G�2w���L�/�RX|j�]O�(P�\]�	�G&D��t��ƠgT�������1$w����~�k����;Z�p!���_���kw���[��잔��}k���w�f"ɬ�#��#9��H�Dw
B��a5������h���b�^�֗A*A�
�Q�u�6��?U�H�}���{�Kb0.3����ҧp>�g51V('�2�;���%(�!�p��y̖�)(��޴�8�VM�Ct!ޣ�>z��71�P���s4"(�!�q�>I����L�/D�vL*r��e�G����X�$<*Ȟ���K�[!)]�i��]d]^��������pϦ�!�.��4��<)�u75&}�I�UU�z�\!-�/�@| C�[���K��G�o 8�dz/��iT^Yy�Yf�c�_�� sZ�‰m��Y���䣹�n�������[�u�)<�5�u@uI���	���� ���xe�/�I/f���[(Z� o��	U�ݙ(0��-h���H8݂:�6Ç9D4�� 6O���e���iM�!�N'�.袿��.��P���f�E�Lg5�51ۧ}p���t�����ɺ����`�D��=�3�bp��+��\�82��Ώ�;��H�`��ur�@���<E\JQ�i�1��,a����t� 䏶�>1�S_�0��-u5��Ě��	
l�78�ٝ%�o��L�\����Ub�t�Ɉ>��7�����$��}��r^^���pa��W��1����<�n݂5�{,�k��C�Y�b|��`����k��<�,u1s���ifQ17��N�:��5�2�jIh�:;�(��G�@�"}ۄ�c>�3!��kw3�dnd���T��f��<k$?I�ĶN�ًW�s���V�>#is?��W@׀�2���ߋ��=ޱv�R����P?���좚HM���- 𱖿�����ݮoH��E)o|F�����ؽ���׽�)�z���].��[�������;15��vS'$T1O�Β��3:�0ق<'�CM�r*��3����h�%�����W�1|��ql@%���0f�j���Z����z�SI�r�c�ܓ׎Fgs4ML�3>�������[�qv,X]��	�.q;rQQ�rH�l��{ꂭ:�"<{�W���N��/���X���5�� @�te�����"�i������AҎC��e�*�W>)�C`��K���Rz%��Fj�c.&��`�=0g��H�KhI-�m��}s0&vB�҇�K���%DĀLϰ��`�r���G�@4���viK�2�=u��l�MY�'�3LK���"�����_kL���e�3F�����t���)2�E�gRT|���1�e�z
�?ean�y�[��|�Y�rV0Ф��^���d*����M+�_jBߴ���,�C������0*�Z��|>&�I�������=S��{�ޙ���A:ۄJFmt��_bR�mF2S�����H�@�����G�?5Fv1�݊j;��P X����qU��G�PX�;��ш�X���ee�;kl�a�0`	�ȩ]���������C�/\���B	T���W-��,�9����5�"~�,�5�`D�P}� e��!<r��h�p�s���11s~��ޖ���T~@��V<�Ji�1�u��31�S�Z�]f��H�N��y�����k"?�]-t\^��Ab���~���S����"^��C�D�U�m'vf< ɨ��L.�2d���k	��?�#�0%���bxw�?qIf��B�E���>��0 r��W	܃2ݤM�cnx^2I�/^M�Q�΢ր�{���X�_F�o�$`�a����[�<���ݴش��ǀ�{U��sA.7�`l��cgw���d���Z�k-;}���9a}��//�m�X��΍lz��j�2�@��4c� !�;N֗�^��-j3'�fw�L�����Q�`avi]�E0��N}<�ڿԗ�v��Ees�$,'�/aaIY�cr�*Аj��5k�*�NJ��I~�_�3���3����+�`W݆���Q.��F� :J��]��.i0��Yju�a��Ğ��i�&j�ʶ��1�s?\�mdȄ��;�n��e.��T��o��>[//�b5�o�5:�w�놷�l$D�2N'�9	6vJ�q�Z4(�cSB�`
���h$Vp�7Bj�39'�����0�+=2����ݧWLZ�DC�yvb=�9�t湆�<g_��I $����i#��Q�`"36�9�\kۥ7�a�S�ũ�iӦ:lY�b!��[�^�g������ ",aN�U��OQ�t�5�<�m�g�?�y�����r�JB�*�l�$��f�Dl���ׁ�y�Iό?^h�Y�^����@��,��=��5"2LJ��F[S�U=�ee�B��K����0���g�N��or�E6� B�UC�?��i�ifʏ��@Ck��H^�;�=����T���]�O>,��J�����
�o��`����R��u���:]�l�J╁g����%A�����@f$^FZ���bh_��%�g5ۋ/��3��|�b���#`;%���ql}4�Ʀh�40���z��w[{�?O���h�
���V�.���i����["]=O�L�,��2��6;�Q�}� �fj�P��P�6 5)���)9`��_a�#0�tX�c,ad��(��&�I���6lK�7����pe6�a���U��i�s[5�Mٻ�e��NNp����Ժ�u�Y'Уbt������I�\Z� /<�(��Czr��N��� ��
��k�2BBp����l��+䒶;������?/}�.�DL��]~�bz@xK6��v~��G���{֫�	�o�׊Du4�Lk��	�x�I1�!g�&�js�X\ud+��˱ѾNX�a1xo��.�X_��D�#$���6(��e�=�����C�"F��я�d0S��$gVH��4_���9�g���ȼ�ec���&��"��Ƌ�-}��k�RG�Z	o�V�Õ�:��	WIK�+�q��q��p�����(UnjE���v�o�y�Yˁ�F�'/k�8G���A��"�<���� d��x��"e�S�Kh��kc���V�,�,߭�i{��Ҝq<�f`y��ߝև������,���
d+�������Pu�|���	��r���Q3��Z���=�d�Cxs{',\�����`��,��ڄ��;0�>v@V���KU�aX	 �����2�+��)��%�Q|*�j��BY\���+��%I�Yx���.�9b���
�J���7U��U��9x��ki_�m��[�^��s��DlJi�M�����xshj?��x;���Cz��Ez�-�����k�	Hט�+a?�� i���N@���q03�pe��p�K?|6R@=?��/�&܅*�dȏ�w��F�����I�LN� �h,���9���@�'ڨ��ؗW��F��:�s'�{�-p�χ�u%=�4s�S�.d~�4�;�lz%�WR������jU�ш��f��R�;ۡP)0�tMU^o�RS	cP}�?C���KS!�a�4�+�i!Y�<�.�"R�"H�t��S)�Ƀ��,E�ƭ���Ј��R�?8 �P��e~�O���O�]���7�<I�����D��R<�c˜p:.���L<�η��X:�a��sEŗ3�H��p���ɽ[\1�t���ʦ�Vc ��8.,p��,8D�ц��������*�WP�e��`Szdڄ��z&H��V2!�i�V�o}�|{:��y�>��w�b��3ǹ-�B��G/�w�>����^��bo굸~f������ڢ
W��w������@v��8��0�e�q�0�������h)��M��{Ԙ6�!��Q�e��|��Pc.d���V��p���X���D������z1�	�(���yy �:@L�<m���O:&�M� @�;��2�&Ϫn�8�Ͼژ�ǿ3o�<�{M��f�N���_�/���,���g�".k*�뵾}�݆�:�������$ ﶓMm�Kzn�uc��=	1�1:PƝ�R��e��P��p�D=�`�uNA��~�U�\�xw$�'b��� �g���T�1ag�m�@��wg����-�(s�J��n����g��5� !Q�+,�jF�V"�y���ķUVR�
��D��\�PR���$���nrI0$��X��Pm:��S{��V�hz�[��~�C6~�w��L�?���N�]��,��靨~�^�v'/r2�K��V,�R�.�l�2f��Hy����k�s�<I�2� �+�ޡ�ӳ��$��6m�GW�<��y$����Y���N�
��1�5��%N�OP�~�a�������T��,k�}�8HC����F0��-��0<TC�7�0�s>���H&�
3K��	�P�;^al8�vD�c����5�ۧ�ϼ���n�Y���RIQ����"�}�Ӯh�$��K�u��OF����^�"�9?8�(:=�������W,�z__dQ�W����l�#�}�H���:�O6�O̄�,�Ī`:g��pj� Ў����Vf���q�n�1��LC��	w(/���ml��[T�y>�/o�]�)]k��X����F0�����N� ��]6�㡖(w-p����A�������y��n҆=��[Q�ȗ�\��ȭ7�������"��_��4
�D)��jjh������&�W���S�7H	��� �T�5��,+����Cxy~Q�v�S%�l����!��;�r%嫚�9�Ջ|O��t����U�.	���T����]��6���RF,���>�a�p���O>D�<&�6I��4����LP�|��fAq��oΧ�W'�˷������8g�@-�*��/΢U�����&�A_�D�1-R��!4�L~AǶ�K��_� �n��4(;~��A��~5�~�+e��^��,���<��}X��ͳ"�}n��|���TX�G�Ҷ'0�\@SJ���Q�l5��0�J���\N���y��`�s0�����>wzHy3���7)D�!��g����6P���=lr�s��nHS���7�����GAț��)&�$&p˞�t|Ӭ��b��S�t�؄�1�X"��4�k=aI,e�����i]��jDG��Y'���Lu�����#�QQ[�l ���
����F����vk�>����A��y�l��/h�����Inr�.���Df^���ȷG�\���Y���g�"�b3��c�T���8�ؾ��_�3w{����í_�t�,�����,�/�^�Tı�ǩW���T=�/�\�qC��\l�;�$����¼��Mw����ɨf,������`��+p�Pb�I��y��� �8�8�����@7#���j_ �`��e�����}#I/.�h~���n��Ԋ+���\��L*>�n6�1�:q����;Y�2FO�pQ�O�$/��C�����IW���7 ��.����,��zC��RL�2�U�ҏ�X�O�cy[>���
������ƥx��6E��A�-��{���w��!�TJ�/� ���#�vM�_�U����J���7���a���rY�அ��Ȥ���i�Ǥ�?����Zn���yUA���r�|
�b��r���A�Dd
�w±}��A�ɵX��CBϖ3�>�өb�]�J`j��mY��b�3�[�ɒ9�>�]����/2�I����@ג�P�D�N.�29����t�\i�)+�v^]:/שm"�G�S|��v�Mf��N�U�ƈ����WR� ^��*�汳��4W亓z٦f�)��߆٩7��B:��I�Y�_��
y(;����S�"�SM�r�50��9'��>�����ru5����&��[�߳A���r5.�Д��y��r#qb�����~}Ԑ.��0'�B��+�1,�84-��K��2�zDKJ�<g��
IҼR���Y#��Ӊ1��g��8��^}�Xi-�v�����klC]�6�Ղ�o�V9s�.��V�|�p�s�-��+� ��ޖ����N)�!q�����&���"�ܙ�C��a9��eV����2�"�$�B��ǘ��,>��=![7f����|S'4����<h�7��ը��u�Q��̙0ה��m=��K�k:}�F5 ����n�!�f;�G�
�뭇���k�1����/x����1�����[�=�C�i�?;��ڍ��nf��HO�7��F���*��W�s1SL��	n���mAgB��%<aP*Pn���]��*&:P,��d��$���� ̉Cˎ��r��w�>3%��n��|����	u]�a�0�)��H!�y��s�嫹�D̩�1޻�8XQV�y>�;�.>Ğz? S��n���v��\�x&��B���]0F@�4b���Յh�Q���ИČ}>�����筓��fL�	r�[��b�O���c�*�J(
7cɘ�[ �������a�/Xs,t0b�8�c���هH�p�sVޱ�O���5�a�b��k9�l�F;�|�Ug�C<�c@�a��7#�q�s���Y�p�Ҽ�]u�HD�">nH��z����s����l7KAc3]�i�2R�r�Wd�M+#�JH�,Dme�SI�Z���r�Ĭ�=IY�U���m�U���v�ȁ������hn|� �B�b6o_*CF�:����9�L~}�w��I
'Jգu��2}�C�Ymʒ�9̣����@��mp�}+����W�d~M�Y�	�4�$��Au7������g�¹�u6��7x����夂�#xӘ�ly�U����4����0Xbմ�M������~�6}Ҽ/�g�i|��e�ug���L���=�9J⃪�6����2�sd��bb�Y�A�w;�IM�'�C�UU��N1�wS�Z�&W�9�zx����<��,��5$N��t�g%̸���F
آ~3�4�&e؊��'��ф�(/���v]сg�� �����������rxy��1Xe�MX~���y�T}�!T�&ýj�������!��_�;o�Ԟjq��~�
&91��ǽ�e���"�/�AM��ڝ}T�Q��'�ʧ�5��}��Բ�]�o0���)H�p[��Tu9��G�-� ̒��7׎'$���HD�-E�n���t҂i��SL�o��܆���c�r8��p�#�x��@��b�u=���\����de(��2'��X��ڻ���(��V*�v>e0���*//ZU���<�	��:�����V�窫��1�)!k})=��3,'������ן�t%fO�2
��^q��Q� 7PŞ@�gf!�T笀P����Iy������\����S?�Vp+؋�yk�u���ڗ�^_H2�9E�V�CbQ�	%�c2�9�����*�#ٞ����F&�:���:쭧���#i�<���n�L;�{��wV�m��u���A�O�U=�ŷ�8����bȅ>��}��Rc�*�P.����#�?v�7q�V7-�/��k�!>�J
�����][�)> y��+��
(4L�<���Ϟ��
�)���@(�!�D)
�4���Q�G%*��xs2��ɯG-�N��R���z��kkLn�������V�J�l�' -�F��%�5�Y�e���9�x$%?����S6X*�'t>4��^��P��Tٽ�{l�F`/v����I���cr^��D�^?��@�a�Z�1���t���| j�0��G�g�8M:O�:ת["@���Xnq4��cr�Zg�h����둃�H�8J~�؎�E0��G,bx[���@���X�)�v#�ZA��x�� ��΢�*�q�����p{ N�Ҳ�XU��I���U+E�e�E�=��KM�X���`�X�Y&�V(�,M#�0��N�Nv�f5��`��P�8�@|������w�/�\�׏���Ys[ŝ9�Ɋ׎�����X�(�;���O�� ���ה��ش,�w����pX��H���.�J��˔�M��?�n-/�G�h�dw�Yj�8�D�����N 6��ۓ�Y��
�,�Z�T�J�P�����s�ǔ��4	u�r/7��,#�W �	��q���cB��~#�ՙLM�+	���Am�G{�N1���5���y.��ތD��m�`�u�W�؅�F"b����۴���yb�9���;���id_�6E�����g�>�N��rޮ��Z�`z26��x�g����2/0Xi����[�H�=b�~b\_~K5Jr�5��f�=��+����{�C��n'��S��(�k�f���yO����&��oz#T��6��usc`�ב���xfk;�pv�\� ��d�֜�����V�'��hV��,mh�N���Ԃ������#���V�Q�M$Q|�`�R�� ���ݯyv�!�����9Ɇ���p	�)����Ex�AnH�>������h�����m���'� G�(N �9�5'�������o��N�k`g	xre7�D�0��\����,Լ�8��%��ƾ�J����6�o���M��2H�7�{�w���,�\��1�Q� 1�Pَ ��MM�ٓ����cc��H�o���؟C�ú�bRl����";zM�jX�����5��D%*�"�VFk�	�ڔy�����j���\�ho]'�<��W�g����oAx)�.�Z��!�e;�K-b�9[�=��.�z(���w�y�'�Z���m��;����XUվ�[�~S6���2r��v�B�"}�ku��(��9&L)�w�UJ�1�{w{~���
�e�B؄���;t��� �.��A�]Ct����f�4]z��ŏf�o�sy=[�����g?�O��ټ�y�k�넰�cȕ\\�pכ1s?�Y�Wմ�ŮB3B�����l�aB�@�v��0@���yt����1J�W��{m��̐���uB��KY7w#�r�?���n��Ʊ����6���]��֕q�RDG����\�Db�:�}��,T8�yva������O�WN��ɚB�N����S�w�P(eS��T��ܩ�9���M�/ݍ�[mA��eK�'��nøX�����c���o�H� t7^����fx_��F�3�)�ϗ�(��.;a��̃����Sm�G	j���9�����' �K�bm=0�� ߖ��z���nmh�vO8���Z
(�����S���*r���D.�
��QA��t��s�D��F�Ug�_�ST�.TUʢ�r� =[�8�5IjIU���R}e���|���HmO�
aaMGaX,9��)~B�[9v�O\VY�?B�Im�|��L��|��'���qs��H�	������֨}=������v��bL�B�c��_,�7Pmq\���N��5@��sSj5��4�:5����5�~��D��qk�B@N鑑�YgD���Rp��VCRjw�/�i �������9P�?��D��Ԅ��t�͹�wz����!�&*��xj����UIּ�����^%��~Q:��RT:����ƕ����Ϋ�4����w;T5+�#�c�1(��A����I�@$-��W
B<��{*�����'�e�u}N�FV� J�e���TY{~���gf:�<w�$m�2 �yO���b�V�5��*������M��\Hk���u.[�ᅝ/U%�p���Z)����BHxb[]�zc�qm�*ދ���˾E�u@ߎzf�C���PK�p���`��ʎ�V�#�>ZE�q
�8	WB-�QJGF<��uX̸̕H{���O����}sa*e��ܐ}0O9R��!͡��m��e��1���x�|snIk�5�!�R��!���a|�h�580{Ά�G�gI��ú�D�.�U���-�BL4�5�����dc7s�;%،�W�QS&�ز�~����+��1��t��{-w�I�����	�:}�<�M����l�n����b�
@�ڸ�����h���E;�b�K�bŭ8ۮ��H�,�w.�y�T���M��.$z�_�IF�W9Bɦ�J~#
JILg��U�9�Y�n��[`y���`\����a�/ N.z����>��Uy�\�M�x� #�rUг򕑃ڴ���Fa?���am3���%�$gSts]���SyޏOB��ƿ�L0��'����sx.P�QLa���>�Q_�t7�))�2����>����cD�wVF�N���è�3ܮ��nxD�6'Q4iڋ�:�./\��q�.�����w��Z��c��_�=%]Q�;�����M4e�r�/0q�]�9P-�rw!� L�.#��^���$�tT���G{CV2�n	��ŭ��լ�o����;;��}rG�ط�]Ҙ����y=Ce=��;��B���nY��[T�I�7�+�.��q^�
Bc(�Z`�[*�"��$���à:�ɞ�O����r�����4�2-��/�����D$������9�O���uJ��M�ӫs�+��$� wy��	T����uR����eN��ply{Dy�[�&js�a$H��j��
�az'��$���s�X��[V��a�(G�в��ݮa���#FZ�p����.������ڤ�'CE	�e��Q�A��Z���4V�0/\�,_)cu��z.��s+�J��Њ���2X��ߏ�LF!�_:��{�{(kV|�)ou�>�ķ�.
�8h7�l����jN�y�iSW�ZO�=%&�@���FhC�`�����[�8�*N�:�5��(�|�1XbZ˭ �8����L/⋠ڋ,Tio��߼q�����0�a \]l�?�4t�p�}��b��Xqb�Va�X�ѝ��J;#���{���c+�=�@����~�2p5����N��g�_�^4�U��v�o�1) c)t#�����"!�����'ނO�Ȑ褪�Ҕ'�NԖlاƕgʢx7?��	jjf��V�w��Tz��Irwh��d%��<��G�t����a��
�Xc��xt+�Fu!`�?��J�N�IB�xL�F���(���{Tu�y�ǣ��b����{�Ȥ-"*^��\�Hέ��yd#�����s��7iV��g�"-:>L�X�/���wMZ��	JǻN�Ac���zڐ������N����"��?Q�h�u��
�c�ux�*� A���Cf��]	U������Y��V-���8��A�~���6�.X�p-X�;�k{�g0V������(�Q��~��(;��g��b���J�MX��c� t�a�,D� 7��iǠ�$ř�Xfl�o���n�L;��5����>��B�&��T�_�69V���ӢGͨ-��5�'�=�9X$\U��
���5M���n�˓)Ӝ���^��p�X�'\C�^�T"$����?��-�;��iυ��t.���դ{*`��#��7� 0�<�}@��=��SI-*Cy��fhH�b��Q9LR�l�H�H��������Jp�օQۼ^:M��}^#���R���D$���!��L�n���i�}�tת�8�T�/gM�Vof�T���[p������1%'v4k�>v�I����O7�
�e��W=R�sֳ��,�2���`�/pD�/? UU��V�h����c��!?]L#�C��JԀR�h� �~�ʧ�0:/=��k��y߀�=�%^B/q�ψޏZ⼴/�ۧ��
x�煹GȽ[jy��Lz���y�99Ͷ7������oU�����@��K[��Qgy �⳶����(h'{y!�h~*�7#�̳$�@7�ΕCyٞ�nh����1�h��6?S�����r@�t(�� "�u�e�C?򬐛� e�Us�*j��1�)x���h<�vj�/�������D,4�Ky��7�\��ض�UVs,l.8�Ln����W%(��{2�;+����Z��6hq����"~_O���̅B���L�U����vvˋ#<I�GU�H��J<��84�'�t���Z$�*��(�(���r�=��F�5I5�P����R�1�����P驍{��	�'xA7y���7G^��2o$���L�t�^ؐ�?�����F����0y��$v��⸑PX��ZM�E�5���qy[7qz�r�y��M[���~����f���Co��;^���D� ���b�f'����:��d{���#����s�g-!��v10�wW�߿�9�'�&c�4	,F2�W�|`���A{���c�|�Ԑ;.�Ē�.+{r�Uj� ���)�wȭ�xr��5ܽ��U`�({��(��$���m����u�����䳱�ۓ:�w�-f_sG���k�{~� ���$�\��Ĩ�a렄%�c�\0]����"�P��%�âDS��Z��CH��%$'�����b��mi��O��[.\'N�	�� n�t>�~�?� I"�7����π�9��.V�
I��|�U=�ħ��܄����5�z 	)s��n��m��8�5g_ƴn5�¶�%�|C-�d@�����G-��_+�X�uE���^�#�O�9�0U��N�����'~�����=��7�f�k�`��KL?�>�n4G]�E�Vϗ�tN��'�}��Z)7�g5, 0#��r�^C��> �"��`�V�M(�T?�f/w0��cP��*c�Mg�:�@s)$-��ƫ�g4}��:�O	�l�g�n]��02�6eL`���0�>��e�..����b��g�g�p����!�yVf�c��Fɳv��Ƶ|�?���)�,����-�ېc�A�g�8�e�Em�4�����{�9 Vg@���|��7?�����g��W� ���6C�P�{0�M������Ѱ6��S\}��ۉ]�>4;ʨN6�6�4��&�Щ7����������bc�km�vdj�3��M]��Ȣ2���7V��bQƓ ������f?Ǒ�|ђ��!��m����ɦ�`�*���	���Dw�; Bk�	�鎯T�o�8��aa"KB�V'.�}�O�j�IXL_.�͖`K�X�KJT���X-�˒�&�<���;�(T�\[qD-3�S��	��
��!'|b��z���v��{�Y"�%��R�e�5�2,;	�r����:�"�E������Je�K�۪e?�A�Y�8���*#�9\L��z7�]!�6 :%�Ebh�:�ȵr�^c���4�l���G�]�h�G��L��QB��odx醊��S
F � ����j�Q�;��_�t��;x��^C�唖��8��O�Q���1*W#��I.�Y�X�nd�`~x��zƼ���;���k��������Y�kc�Th&���I����������.摱_YƂ�j�*���$s>�k�>���/�%���#~љ,	� �(��F�d�A���lƵ�.ve"��F`��:8��-�S���12��.�>gR����ǣ⌿*�e�C�A�N:���<(�׽�����\�yj{w����o BrYݼ�����&i���`8Y��98��j(���F�"�4��[��S��O:���*�q-��lqUg��%�+'`�/U�
�q�膡��ώ�&����w�|��y�7�Tɓ@B�e��򓢕E�Ą�\j&5s\L�$_w"��v�FM}��s���ɱh!�F�Q�8of��I�����@��s�����[:ڬ$}�yTtR�01D<Д��k[zp���cr� &����0������h	�Z�z��/����F�ڹ>��^����Qxj<f�X!��*IG�Y���j�?��p��P3\7�� ���J�bߞ�b��6��Y�w��,�웂?.�l���ߗ�	��� ��y"�}�L�D��uv�ϻ3�v�L��K��t�R<�� 1��S��b_�ܨ��Rp��1�u
[�43>���l`r�錏Н�Cx:�^�0N0>PU�QN�,�s����$t�*rC
&>A��A<E��3�4P��.C�Z���m����R�����(nc�P(�K�3Hs!�S6��匽{�Q�M�-����9�#�iқ1��2X-���@AL���YD���⳹�$S��p�af�ч��$�R��'�Π��[�SkSH��}���)O6V��^p�� k�-�N��qוJy>�`Ȇ��}�GpYJ�����΀�x��:V����`����.[w���ϋ��sd8�\o�~Mg8�O�Ztu�~oQZ[�Ҥ-��Jq���'�����
��PK��df�2�E�U�[U;����́7�*��u�C ���#��� ��}��Kmk�3�;��h��pm��n�����By�Kk� ���LgB�'��RE�4�[���6%�&n�'V��\��*��]7�9��6'��^4�S�5E��]������*4��Q/�tO�&��k^�uJ���n7sr9��GDհ9M o:%wyzᠭ�-a�j�y��ڳ(��L��J��
�`�j)�.���}�M�k�`�kd�55X�ŬTj嬸4p��
ͰY+t�Qn�ǫ%���>��2�ZR�	 #fr�t�1���e�?_X��k��-�t�F�y?N.�	q�aQ鯞�L���ǘ����G�T[s��q��c�	�u:��@B*�_F?$j�Ң����B��c}�������.�JλQ!��_�-uz[�f���Ƌ�o7�5��d&�"'/�(�v.{�x6�Y��zV�)��FVy��Ne	�w��t9�7���_F�y��R]�b�ϙ�K8"IGJ��NX��X�O�d�;v���g����ܠ��kp���/�{�e�5���C)9���
����|� ��!�T���֩wI����
ziK]�~��sqQXh�/|��K��d�zԙ���dc䌅(�iۖ�3o���
G���Uhc��<{�p *mLA{WoI��睤�0�u��=��9R����
�}�",��eb�����S�����ɏ���m��4��2��������(�=G�dF:h/!��ή<+"3N��1����"�m��i���c�Ӫܬ��9N�,9�B���N��V����䐅4����O�$��p�"�f��OE~=�bh<d�S�;�>���Rx&�ںki�q�����V��� ?�W�x��Os���k�@�K��c�`�����}|�\���3�S�f`��ҙ�~���Y:%6`lq^�)l_2r�k	�	lP4��k;�MQ�V��`G��w��i.1t�N���D����Ӯ���x�0�wo��jZ��ԩ|��1`uR���ٛ��}�,��V_5��e��d�C�A&۞w�ߺ�O���6�H��V�Il�V���>3̓$�������-k�#��n���?�6&bReظW��ވ��8��K�,�Cn�|��W(ܣW#Ԧ��T�ic�l@��bN� `o�O�z;GI
;8�5���� 4�ʌu��Y�LRq��!�B�%��*9��'ǁ�ͺ�ޖ��'�g [��E����n��ɡąT��c��B;��_7AR*k���Ja���q���Om2K�������#�=�H`:�g���s6�/\^9'&J�
�qL�SDn} K���R�;��������}�t��N��Ð��$ҧ��MQ��_# 
�>�7X�~����S}��%�Fq�+�WO���22=	�$Hbڳ���F���~�����!��3�}�܅l��C��Ii
�O���]Jj8�T�:��]������G��QzHP+)� �9��I� _�B�7��)�i���T�G]V\��Fι<���
��giX�ߐy�T��JF6{)�$n����Ι�W�Ii|�{�:�fg����{$۫eK'?��D�쵹�g��h�&x?��0 ����s��=�5'�?�h7"��ŋA�����~���~�%�0��>]K���2p���8���n�k++��{�V'9{�4�q2�Υ���x[��b.�FS�ƎM����l��&ހ��ÄK�E2/�b�6OQ�vb�kηsqwٜ�Ap:n�/Q�4�x�a�\3����X�o��,���E��N-��R��23�FK��8�����`8�!�ҋ�4j0���"Gp}�&������d��G�R�hA&pk�L7W�M���{�9�2v�l�Bʱ7cM�v[v^��Ġї�C��fdĠ��b�gר�d=�HC�ԋ�t�3���u�ܻ�,���$��8~��Y�Y�N']���D�鄡�W���m=���Ў���1�*�5Z�)l���M�Р�P��&�;WE�z�#��Bg*��խ,���t��������Nz����'�j�~�))g�ҫe:�㑦�^��띻c"����yFO+���6�ɍz���M�@�~\����7���F^;~�����:�w���Rҥ5e���J0�C(U[���t9�=ri�0"-���;ǟ>��W��w��kD�+�������^mփ����h��}1��~50�J�_D�i��l6�GMI����L�cH�=�ƺ�Dn�=�d\D�[_�K1}~��݆$�=����x���_/�qwӽ�,�QPöIͺ�����/x���[�?ˀn8��v|�m��f�h1�⪛"r��NiB���{D�,��^T�A6巳��L|n;l"�5Ѵ|�L�:�_v�$�"t�[�dS2rVw49�T�"���x;���z��$��sw ��6Ԓ@wܮ�""~�:��s�S��9#Sηw�k�)ĳ D�v{5H5�!��S�|�xU���X��&|2���xJ�p�����aO�A�nJ��d�&�x�2�����OJ��ΪЉ���C��
h� uS|��Տ��tD�!�N߰U�燦'u�0��HyZT�tV�'�AE���j��j������27{�Tؙx������ޅ*:S��6rqGN����ş����G��sS���������}�^S����tń�Ȳ�?'m�c�&��*���y���8<WzFT��č�Ĉ[�̎	�zՒ���4˅~��5�/��"�٦�] $�8�5*����}�ڊ�����IN�z�/��j W㫺4��<(�R��=�����- �Q�`�{x��2�-��N��b�=[#uT<a�P�$�NQ͊�JJ�sVf�\Y�����[��cNА��eߋ�Sm������jlFݨ�UҝW(�V4��Һ���"%j,\+��g���F���� L�B)��+'�ck�k�\����O�cNJ���#e�4��
�:z�'�y�	�hΘD�
��c���s��sn����[4A o�%���w��ݪ�aD��J?�!akuӾ8�6�.�J���`��0��~��IK�MGѲ�ã��R��c�� )tA�`S\�Q+k'"S�����z�3ԡ�4�ܐFiÕ�"^DG k���%*��$�pE��m~�G�O A�Y���U{��6:��	˒;G;�шCR�d5M�"�LJuL�V�v#SI���w�	��m��薯!W�,d(:U�H7�q�����J���_��\nb�'��K�Z~��Gv�y*J��&[���E4ԙ�aa��j[ߔ�J��ؽ�f�7�zv΁Ș��OBM��k�\NCEz��#w]Ë?�2�B���=�aᦈ��=eo��8��e:S\߇[�a�ra��'��> 	�#0��	#���CZ�����2#<�@+h�LZ��]�"�ZQ��0����%�Q>��6y�"N��{��J��G��r�r�{ݴ|����������QSBA	�2�g�̄�r�U���P�!׿����.A}�SסQ�\�f��N�=f���p!���D������-D7t���V�a,�xI���y@�@�mx#���q��'x��S���T;Z5Iն�m��!��nSRN��emOwZ4�R	�W��=��&A�C�f������g"m�E�ڬ<�@��k6�38zѠFX.�#B��}���� ?+ohi�Y��pUK����'���#B���j.�v�x���h50i��I~y�1pjS$p��B�! r��������iR������T+���+���Y����1Vpc<P9�>��'���(2��0�H&I^܉���mo�����d���\�N9AD��P�6�s�a�-u�(�h�<�l���H����_1yI �*\`,Gո\�j�>�`y�>�=��>©*R���~sN.�N�.�Pc�&�Q(���r�TJf�u���g�:]׍� V~U����73ܐQ�`�^.�vW]c�
u�{a씃v�B,�Cg[���&cY#�fH`�f���ݫ��,ˢ�����.�@9�d$D�f�rv�Gd�_3]�w�qӓ�w( F]L�J��ʑ����Ôt �G�R���*��㗼?-�cV���U��U��<앋�Y6��������:�ɋ�b�{�QT0��
�|Lм��6(T���jY�(���v�3�;)�3�9w��{s�'��!��i��VG՗���_�'O�aWP`���uF]a���&��H����s��Yv�^G9�b�3��G�.K�h��%	��S�2/Fz�!�ׯ��Nұ��9T��B�KF�j�@�O�&Ƈ�;ZW���'����`ޕ�5�=���TqD�s,���WZ!��;k4�l4�3�������{3#ۯ���E{�X��ta�4�{f�3�r�� u���4����6�G���6�LT�#�9�n��o>��AhU2�غ^�-J��jRCI'��<p]t{LdR���
�u^�s�J\�Ɛi�N���I�����j)F��-����20I���	� � >��l��� �,dV��~ua�N�gU����n�ݶ�����+|����r|��p�!LS[%��bw�san��Ib��J[�BQ���{�i�(ڌA q�����l�����J��gq-b��,���	t����b>�j���4�j���?�\P.�'E/ߤ��7mV�Lа�k�9�;4�s��o'��p�/s�v����Ƀ���� �Ȑ+G�pM�7�D�3x"��t5^�S� q�R{1��W�y)�a�Y9݇N��m.���C�E(X�j�4Z'w&M�SdX*�tN���kG�+t����}@��uY�����<�^A}_e�]�r��.�v�s�9��F����s�Pc[Z;�C�=��:;:����7,2V�P�p�_a\/5І�O�{�jRj�e��p�Kd���u�Y���?��0�ʀ�;���Q��5jW2[�_�˓ֹ���{�&�9`7����f#�1��v���Q;���C�_�rM�h�߭ ^���C������t8EDk�!dE��杸�/yb�#3�����6�	��h�1g���p�u�����9:��T��R����m�!�"���aL�#)�W��yE��΁�=�	M�_}R��LT�H��u��Î�G9.���{Ks�0TT9w�s�]�N����F�["���=|dfu�Y���0���黣!:�(Y��k7'� F�~��7���2|��L,�B��LQ�J�ɞ_���J]2g����!~�Z����T!���@�^��J�na��k���#U|���Y�����A�2����%��LF;I���A8l���ز:D{�m�KT�	ȴ���\��]sٝ=����>�*�;s�@F����\��R��i;
�J-��?��䗁2f�-
lqi�`���C��+���s��_(����!C+y8?��lr�t�k3�}b�=����|y+V��2x��ґ���m{���(���˾+�*=��nT�p���o���uϚ�V�}H���5�>P��'r�v���-8`��/~%�`_4����ݚ�@������o����-?�T�I�'�d��M��0ty�k�@ȉl0����5�r�r�5fR�J뫀��D&�E�ԛ��VFLr���r�z ��K�u�&6F"�R���{Wd��S�!�К�w�Z��L(L�<����zdh�]_s.��YP��M�2=OtR�(f2q��%a6|���E��&��2��C+�|jk����9��� N9Ѥ��~�AW�C�rj��H�|��و�sɼi����g-B�34{�$�6&h_����ѥ{N5Jy��a�c�6�)\��ft�Je�g��?�k�",CľQL���0,	{�ϿWE(�荍9��r���c�(N|�x�������(��p��ڎ���r��p2g�V�L������4�*4əE�s�4C½V�R�P��Q�X��&�k�VQ�⾃�$ck�Bi��`���ItH���~��j�j����X4DWo����vn_ܦ�0�Y��胇�2
���g��V�3"O��Ddj_j-8�l����x��BC�6��5�����۟jG��S�ꠅj�m�%��=	����X����Z4vW
7+�%��M�2.�AZ��I˚��Dʙ�,9�`M��z�G7�
�8���g6�ZH��Ⱥ�X��J�.	������m��/H�B]])VfS�dt�(�Z�Ndց�s�BX���*#���Xv�u��N�bj���6cۘ �侀,�TfYp���qU��W��㸽z�^����mD���`�}�c�v���sY�4���ey|S�
\6c�_�����c�Ŷ]f�&5 *%9H�W���4��,R��% �%^"ǅ��"n�Jj�W���̃��[���/C��QBg�������)��V��t�H'۰��X�G�)�#\������Y9��V�o��+�������s�M�l��Q&��9�%A�q�+��ř2E���%\п�yh����*�q��s���S�l�����!�ABx�(��q���dL}��8PAp��X�U#���^�kJ�4���	%���j��e�� �fڿ}�.�INZDM������� �E�/����xeO��KSr0���U{�\�����%zJ!	J�±{�I9�T8�.l��m��c3]Ç���$�B���y���O�@\#c*s����yN�fs�&��~^�S>��L�]�v��c.�9�V�'cD��M���ps-��}�VN<���(� TH�If�>�9c�j51�	�lu��i@�����9kE��H���j
��g��T���N�&�[a�SQ��|Z�^s�<CO�>���j$pP=w/�lGD5��w>cl[L�T�ϴ*�s ���fj�ۙ�r���#2��E�ӊD�;Yo��I���#Bcﾚcv�����`�Xd��%��1p������z3y�D�1�~e��|�u�x?X�uO�����7�ge�#x��N/M4�/-�
�5���I��l�O~�	Usoi�!��Q�t��� .���p�Jr0r��|��{!+�?�J��_B�c�����c��k>����#6�n��}g/�&�.^,٦��]���p�.�CI���;���t�V���l����T*uI����D��S��w��v���T�$��]���o��U�g����ay���R��ڿ���W��y��pT�����N�O?�R�o�����<�v�ɬc#���Y��$��Ɛ� ��Ϯ��i���Pǒ�����|�Øb�����,��e���������L�b����״�Q�೟�s蠟y���6��	x�	�\-���y����y8�ėx�U~v@2�-����ޖ]d�Y��/�۔;�-FY�B��w¶B3���@���b��HAg{���v%�t>H_�>��#���}�� 6٨~���i�Xr��E���s���վ�m��p�|��7��}è���\
ύa�:��R@�X�]]S�){]�V�w$Mbu�<�t!6󢘝�et����;D�=<�
/�1�2�y����љ��
�G�)��s�ݩ>�^J�d���d�V�G���OI.�
:a�n�� Z�We"���(I6��g�.��5&�l�ҼFR�EǊ��������\܆���KW�O	c���4m��Lg�21��oJ�͊ɚܪ;�����ػA-%�Hk��v[�^"��Z.���R�������r8�!�/��L�q��S%dk���k�@Z{������h��B������F�K��#(]�(��D�Zϥ�(eǟ�N ���+5 ��e3xS�r�Aլ�=���|����(8x���ΰ�#���z]���x�D��~Au��>8T�X��� p����� @�|�?�0�Z�K�Z	��ۊ���Ӻ��U�^��p IJ����oAh�K^O%����=��B1�Hfjnxikx���Yo���3�� 7;LTi(g|�s���@��DrA	)�
<M�dy�8�p�����>�֖�m�������Y�]#�Pz`'�� ��`.�޸1b��	Yz�gX���W���bT	V��(K���_K�U:}�^����1�;�I���ꐣ��J׹�mi`�.Q�[�����2Hp��T�}߼7�
M�"�}��NK�2o"�X�%���q�p�	#-��`�id����2瘲;�Q� ��<����+޷�S���ٺ������d���w<��g��*��H�`��4\"VlP��dJ'���4	�+���F�\�����`{�zs\&mp����f�N�1~��ޞ;���#Vār�<�f<ap
��"�������暳z@�Q�%D��p��e�q�z�������l4�AH�#�e@�⸩ӥ3�(�y�H�S��ы��&����y��^l���}+��d�!�a;�=|�e|����B;�+��e���%�ۍ���o�7��e)?��G|�����ٿ)���t�W���A}�t;٪�� N�����KK����iR���y�Ȫ��I�>���du0�A�!m�SA�M���6���a��ה+PzE"�o$�x����ϭ�b���������)c�$�i�|��d�~��	g�/ex������UBW�x�f8���u:� 鲎p*�� J�!��n�����6\QL�U&MA ?�I1�PܹP��T��Zވ��M��{K�)AN�Xj��u�ܫ����^���`�p|�����0��� �|�ev9d���cep��u��X��iT���x�j��eű�1�0��]�۫�94?na�t�H���{��۹��s�hǋS�f�ВR3[�����6�,n�I�@�;bkh���6��艹���L�ч>Е}����9(?���g������)à�@[E���8c�sS�DTQ��N��"�$�
Hs�븀�I�r.=���YV�~�60wu9ql2$ڕ��M�t��9�������َW�(� m��bA����hX�hd�#>l�����m_�Ph~���v���s6��2�x�)�GO���Ϧ�|t��BKq�"�
�\Q Ĵ�j��g��ŵ��epꒄw��"����;2ly[�!��uv�vl)T�u�f�&0S���hw���*47>��M
5���x��:�(�]��ac�[�b'd��ȯ�7����y��v�7M��gФ]d�iQ��]"YH�J�E~���ĸ�ɘ�7��z5Q�FJzjv;g�T4Q�]��6���|5�& @>'���Y�49����A'���Q�T���I>aR4�� (�̄�G~a8��!F��S�#ix��9L�mҹ�M�z��ޥ�ik~���v�tW�W����a��%ީR�y��6�d���0׭Jm͝��o�Cyj�)���Rq�`�*�$�Ue��X]fC1��z��|>��=��=���D�b畊���R��%��v�s��_6��Z���Ls}.t�%��۶ݜ�W�����\�\Rc�LؽM|�M��؁� $7��q�:��n�n�w�UN��ѱ�U�)�,�����'��^���!���V�mQPz��Ɔ�Z�̔a���@�Ā3$(�H$�`\__s{�;�3���ہ�b��K�>b��H���[�z��7��[0)���l�t��y 8A������C��@��NEo��&i�m"�aig�w��i��c��+p�]�J��&|}�˝�i����g�W�h�*��t�K�W��F�����U���k�}臡+tݿg��o�mW3|d()��s�5X�Z+5�ٞ�D|�դ���8 ��U�n�h�O���u@P���$+c����W!S`�T*>T�"3�ff!ڥ�l2� H�<��2��Ϊua(@��c�g~��&,V�'(�A���f��1�9�!�gy�OG48<��mr|Lo֭�8�-BG=2�a��%D��N������jS�Rv,���2(d�$z	�`��ޖ(Dv�o���(��EZ�r���C��B<�w�� ��r=4�J�%��F��H��x�t�X}��8RTj���4�!P1%�dv2?���WD�	��n����GHAT�>N��ƻ���(�PL����pD#���|�?��� �P0F�Y��t_����W�j��&~��o٧����DKJp_�����%4�w9s���Y^�3�48������H[-�����K�(s�� �����Ŵl=���{��ޅP��Ib�DB$̒��]qr�,a���u�_�� ׾zF��Y��=l����	���g��<?��s�3e��xQ�vH%��0���1��d�Hu��-C�~4А�����O7��vu��QJ���c�7k�}���8��{��b�a��"Q�%��������Pӳ�9����{��B ���W!uLK4t_M-�<�BT�QX�Y��ȅ������D%a�!$e��ۛ�3�]�ȳ�^!��8�O��FN�A�?,�&C������m��F-��n�@�hjp��:������`���&+�P���oQ�~�Ȗusr�iZ'��y�������?#����LJr�(����\��y�{�Y G�K99�>hƵ��{%��FE�������S:�I����C��5�6�[,I 
�pӈU\��;����0�J����y��^?�>�	��=��8a�
G�5�^��;*�xDWĥ�Di��8��i�v�3M�7?�+�a~z�0(���gJ�$�ج�!βteX��g��n�5�/B,"�
x�WҤ��r��nHZ�_6�mkG'"\3�9�C�=��c�5�))�[����o~��nd ��F6 ��0��Z���ya����	
F��ݏx��*��W�~_ [���K�iƝ=�$	���b���2���f�u�L�ЭB����`,0��͐�Z9얊��{�T0�&��C�+}zt"�؏�w/|��֒��>��8��� ��S#�H�u�c���eŸыDc���:g&���9a~9iB�"fM��
[�2O�M`�=V�������2���D��q�=�v�e#R>��w��+B����3o5�*¬e�c�21�f˓#R��R�����u���H�6���H����ֳu�pf�!<, t�M��J����&����o"�,� x<��`/f��ө��$t'��DG/G�3���kN缜�Y���lJn~sT����ŗֽ�B��T�4r9�k�������;%#��e�K���Ul�	�4��*��!�-��>�7ӥe����ϵݥ���7�1����[���O\Є�'��� cXfD��&���P� �aT�/�XP�gVt��/;7��	_G�9���V�L$���4�u�ز�C`�jӫ�!
mļ�ƃf��kx�g��Ig���͔I �z2�!k����'A%}O`�R��zt�zI��:Mi�k�"Ƈ����'Y�|��
7��
'X��-��0����.�%����KP���6v,
�d[�3� �<pUI���#Ƌ�j*&����Tl�\�����q"!�Eb��$!�/�!rx���L�a)��F����+��a����uE"�)hd�F�:<�k��g�`9�cCY�?e�/~ꞁ����	���`��o�j�� ��������vD�'�H.Du�BfS>j�,&"�2���O�]�>�Ϣ$�T�W��L���r��e�����[���χ�(�zM��b�r��{K�U={l�O�m�r,���YمU9��3��m�=0ME�FaStݑ�P�i)�,��� �%�f��]��ɝӋ�g�gf�d�mj�?�A�%x�N���T��l+�?V��A�_��?����a�'j�8,/�,A��N�������j��ƯU܉ե~��5��^����������<;�a�+HX�3��cc��2+��P�S"�d�gk0�(,�=�շ*�`�q�tM�a�V�W\��+u�W�^8v����I�gJE���&j���j3t�(���
j��6�Zԝ�(�@�dԟ��z����a������q'�q-���v���KJĻ0j���
{�[AO�&��a��@&C�Ԡ��p5������A՘J昸 j=$hѬ`f�v�LΉ�	�Se��1@���T�>JS�<���ȚAS�Uۋk]��=K�Cd����� ~2��{�"o������1�nInm�Uo6�DA�\5R���H���4o���� �;�+B���
�ǔ?c9q��g����}��X�5�Mb�IŊ	9��ç��{�*��._k�<|�t�FR��sK�����	6���y���\� ���׀s�Y��9��Pb��̤7���(>!�V��LQ�9j��^]9
�����F�v��Do=�f�k�bT�.1.?���!2<�ピ�w[���( �6z�xq�r�J4�k���管|=Ѯ�l�T酟�xH�
ˇ?�"<�6�_ǰ��uA�r�<��Qn�� �������J��n�ɋ_���1>�?|۵��S�ӌq�Ǭ��3����(߉W��&ی�Q�?��s
H9�6� �D��VMҎ����a��<��$��*�$^��u�+�J˅*��y�x�H��� ���U"O�M1Y70C,�YT�N�:�]y�-�{�4f �C����7�<g�h����۸�@4L`������^W�B���g|І!�Ĭl�D{��[�M��c���E���MO�>���1���`����%�0��ёp�Sf�-,v��|��&��0�K����-&1㟢;dYC9Z��І*�f�<7r�����я3�:qRE�l5��;�Uja�Ie�ۻ�v�Y>qȻ)i�%�N����/9��܃3Z�7�r߯�6E\u�B���V]䭐Y��g��j3��(��5�|�98^��9���?a��2�h0C%��9m�43�BUS)3&�zy�mkm���5�,����樀��X~�(�|l�z)��
�Z>�����K�^����w�j�8���5���ZI�E�3R.�%iKh�嬮�R?���/��?G�42&FϨ��`�  �y((�|�ƣ��w
�g�!Դ]0�u����4�ց��'����+�t���'��J㋾uߐN�RΠh��}!�	�������WyZ��t���WWAan���/A㰘�y�������x��6*����R������ȢK�Q�X��S�<����<mV�%��S7�#���5�h�'|etꀷ�����p�td�y\��c�y|���̵�ML�@���b'���5�[VV�,C	�(}��{���\B�+T]X�V���p�������: in��!�@[u xuC�pm�����:W�+q�Q�) �������,01�T�~��txm�r/�o���/\�ki�[c�-*@��!��4.@-ṵ̋�S��?u�����"2��'���:���g�+H�F���8�a��p��1I����S���"��~Һ�4���F��� ��W�j^V��``��Ԭz��p�%C=���|�����O}�n�̼(�a7ạ��2a��Z�����S;��a� J�>�Kgrz^�qR,�`6<�g5��yx�b-y�=P�~ʓ2���vXN�A�D�NW���D�h��0���CS"u��H�.k5G܋�T���:ڿ�4���e+��<���5��."�b'ݽ/�Ɔ����E�n+�Ԧ뭬�ཾ���'��bZ���cz��gt.�m�*W!Ӛ�D���|p���r�V�����B�0�7M0�3�}��(����-6���k�$HE >6Z��q�K��xr_An�A�5�2 �e��L�O韝��Apʈ�v��8��tD�.2�x��X�{�Ԃ�Ԭ�X8�U-_JJQ}�W�����^�W}�r���"6.1��tDDny��>�>^�,/�h�����W�i��w��Q7�]KN�wvVB��Q��7�H������h*���=�hD��>ny
�w�P��#=��M���#��.U]�|đ�RD}ʑl�t,���hQ�ϟ����!�h�g��ڨ&��vk/��T��5���]�GR15z@��R�����$@�`%�@�0����Y��7���Yv���Y�=7�{�(���{<��8K�/3������Z&S8o�&z����Fv�
�u���;Z��Ś1)ʝ��>f'i��}��p��r('�1�K�;�X�k&l����������������E9��(��Y�/��l���*Hm�=*���{k�^d1�g���T?�.#�=f�Ҕ�/�7�@�|/�o���1�>/&��I��̊ː7ts	tv׉���ԥ�YS��5�
	 8C@T��]w9w6d�������7�]f�5�f�f��!�������>W�q���a��ܸv�Jϣ݁ F�\!V�֬Ƶ;����=��7*�Q�r��x w�UC�~�f䍻�2ɌW�O��^oED�3>q��Ȫ�����~isG)	u$��LY��A��<옩s����4������Bx�~ۍ�󆑱4���L�2i"��� P9��'!�Wd	�S@�4��p-,�:!	޷��}���d��������՛��;O	-�����n�p°��u�o�r$�8ߡ���75�n��qɪt$��5w�E�7�x/u�('G��i��T�0�?��ӽ<�"B�:�o�N��5�}k�wO@����?��~<$v'aK˚Qnqkr�L7���Ὃ��LH�n]�@��$���+5no5;�>T����B�z���B< ~Ǝ0�A�(Ď�GYX����gts�m�V��`�K�Sɀ�K��f���_�����$���ɬ�1�.��eD����Fv9e��y�����qCA�l�k)5��hj\�@E�E�[κ��pe�b��;���:2w��m���a�6�:>.���jB������B� Mǭ/(��x����Qȡ�z����C�͇�<������w���V�8����ʑgi{	�]��7u'9
��0Ԡ�H����Ok�にC}��izIS��%�H��u��n�ۗ�]e~��3櫃�\7e��R��:<�J|�zb(2	� ^H���i���ip�;X�έe��L'#�o����BG ��{I��k��۸��4\2��[19dc:�2Q|�ՠ�pچsz��T���ފ����o��ܡ���G��c�Cu��s�0��Z�hB��IW+|�+﫳��
�
6�;N�; ��o�:u��R����"����6T�uG��qR1��Pq8g�O����'y���������K`� �(@�_p�����M��+�ѵX����9_m3K���9�/z�`��9�mq�j�-���3���iة-�OūY/�pC#�����K�]�S.�[��'��ÜӪ����
f�+�u�0���:j�`�D,U�G����z˯+�ܠ�Ur�Q��\Y{/���R��>���Fl�{�&�Y觯�0/&��gu�I�t	�n��hOo ����O,�K)�=a��2�,���@S���o$2��oZ2�)���dCG���3+�'�8hc�\�?��=�L���Z���S����D�O����޲ؽ[��+��|���Q ݡx��TEqar�~��F��k�m���MSJ����u
_5(�TY�zY�Ȃ��A�v��f�dcÿ*l�&�9l��>9�&�Y˞F�`��i8�r��P2���͇#{�H.�Z��# ��uL)�gB�����4��`�R:�XĜB�^].� d�ǍX��3���)�����Wq-S����������L��l"�X� ���{*_�����`��2˼��Z��A�h�����p4.�?b���s�����'�rST5�,Ă�.2�+D�
��f�N�'}��.eH�s+�b�R�f26u���4N���-2E���Jηٮ�V̷�۽>�sNh����$��gύ�,V��b���r�^p3M'�7���a�p��<p4�:�O�x���1
��[����Io�l�d-��%2�3\̇6����bl4���]c�ֳ=�g������͞<��ݔBۇV�ӉLC)X��60ˆ;��_�Q�a *w�Ӈ��Ѿx�1< $�U���s]���kwHc��� Ƹ�W��;p(��Tf��q�o�^IVd��`�AZ �pywH�^X��������a2�OJ��`����3�������i��ܐtsC��� ����r0�Jԍ�(��#H�8`8��;�/�tπ!/�}BA5K��/����c�a�n, {euU�冧�!�95����GΑ��R��ZZ��:�i��C���,D��ס]�i�-�QΌl���?e�N��W����_Y��㼩���I���w	YC�!~!���1Q��jY���c�F��*�$v�iA������ai��Λ�O1����gy㋰LqG������z��Gi3�1 	͌��{t�����Uυ�1R�E$���Y�<����#���h+���E�ϑ/h�m,a�ֲ�'�����F4e#Ʉ 𕣊0��>��������8��5�|lQ�	i�N�ޱɲ'�-�iN:��UT3V0��~/��C�9�'1�`����)n���9��/�0It�r��C`	�����T��z�u+'%�`%u�	�ʙɞO��N�'"�35�*��d�P5:�G�'�bcr�5�6�_O���=b�и��:�`����4��O-�㑺�~���5z�n��S}U���pI+}��x<�s�v,�J���O	qW���wY̦d��@�V�թ9�t��ė'$L	�u�����ӂ�ӵ�T  ��HN�E ���4��3k"�������Qm�#��t��:#�}��I�A�!:K�A�aт�jL7��0�wUAY���M$�_D����U�v����Z�u����5z��_7�HLv;��G�Q�I�<c�Ґ�ET��!l�qaB�3����,b��*�~r�����0}�_)f0h0@���f�n�N�����Zv��?K���prv%d-�R�=�G/�C��y�dh
(Q�7�P[x>?�ûv�|W�1߳)��}+}A�����dɺ�Җ�:��������%���8���4*8fqT��썉{�`�t��[L$
Pp����)��<5?G ��"���G�z�5)��ngq��=��d�pY����1'�����m~]�/8�1�:�f�z�[�Kc��ޢ�����&?S1�9s��n/ѐ��S�'�9���^���p	�A����ac��p���r��I�h�/{��Q�:)α���A&]�+�[�z g�>~�#�▪��u5�Q ��N��<���&��?���^1������������P��~�w�G��y����+���M�aѨ�p7up均�<��|[�'{W(\~�}�T޸�89mrݸ�[U7�ޠE�˝�~�y�4��'J0�*5��SE��ȸS%I����1b�L�˧ފ^���*�~%�>E'�0��]NN���j�3�{�Ӫ��ƃ��]wr׽|N�6���fs��AO��+�7�����l��,��R*[�ؽ�ǭ�>�%�*yY9���Yh�$�����Zj����O����t��)0< ��.��cơ�MT  ���b7p8�$�bv�i�d!�7�$�N��D4ɖ�J���**��}9L���1�����E���2A����b��t1:��õT̒��xFZ	q.Z��3	g�	�� ��sU�tG�[�М:h$7�T;�;�C̃Y�N�������@�/$P���pT��y��;�v�<��hE��2È�Ł��xX�e�W��|�FҔ���C	��\=��Z�N{PI>�ЩN������[{��I;�qo7��d�ءS��|HaER<ֶ�X��c^@w2���sA۞*q.��+#�l�>/Z�!|~ȟ���4e�ncٵ��zI�B��?���L��ɐF�--.����U;/�GPu����ż\�IL��}�v�3��DK��W���������t���j�-�z�!�XA �TTY)�ꁊ��R\m��}$G���n���]
�����/6G�aI��ܱ͉�,
�R12]0G6e������,+"	�E��=,򙯾�J&�2Z���oF���<9#0Jb��E6�+�����ސ���m��5�a	>�]�D�ؕ���Hkfڌ�?�ä�W����\�vf�w�d"�(��7;$��M3Zl���>�{Zg����z"=���Za}���'IE��~��>�ǫ`H�1����T�OV����t8�{��*�l�D��Q-�A�䓼��& �U�4Օ�%�l��Q>NdK�A�K)�[����S�rpQ��ۘ�y���F-�ni��w�	��y�&ZU�n?V-���|�󻞝��>֓��S�u!��-��R�A�cIpPߥZˬ��#ߞQ�;4RN��u�^�H���N��u�C�3��y7�j������kD��i�k'����t�Ģ�yN�T�1��V]�w���٢��� �*�2�i�p���6�'��g�4K��	��a�#�Sگ��$A������c�Y0Uެ�ѝ·���w��ߖ���Ta.�s�8`ԣ@�-p��h���̦��~ ���(���}Q���Z��U�j�y�gs�)ȃ���x��Ό�9949d��5n��%漕�i�e�_�bB��~�}�T��춉�jfry�'�Fw8��c�G?��\�A🠙���b͞s�wB�C�i��}(�ß~sG�q��Y�c�xj��s�
}ǱQ�^E�}�nj���PI�=s39P���Q4yT��$[l�w�3� 2��	F��V��]hٽ���txb���.~���}�z�^s3�ڣ��h�&��f��<��	P�d��+�%�nd�Ś�U9�g�xZ�m�7%�e$5o�3���#XP:'z}/c�,�ɿON�
qa$E�����Y�k�gR�G�����$��H\5'd_�3e��Ubq�R��k0vv?01�T��ȋ	;)�T<�W2��A�&�`Әu�~v���ENtt�>Ll���f1��_ĺқH+6�OD�|T�������7?LM��̉��pW��=���*�n���j�.�8��ښ���_��"˶� �mZ@�bd�D"�V¨[�̪�UW%�E8m �d�_?1�N��
�}�~ﺃ��l0��NC}�g�+�X�`?=iE���F>Ҕ�P�yv�u?����s�i�/І�s�/��4|\�n�
�̭]�~�Tİ_\6�?��7�*+ڠO�ɠ�7	��W<3��ٗ�ۺ|��e͐�A��Ėk�|�|�j��r�4A�p)�Z���p�b�V���tJ_�MI)���+ɓ�c&��r�h�"�,0 ��=5WoR�`)xS��
�6����u�1�Q))�,P����]$j9_�F��h賛����`��
䳝���n������Dй���2/|��X"@D�_������2{.�/�t��� f.�}�/��S�=��?��p��G�q>Fp-Vp�,:"NUc�H�J!��F����lGB�c~�I��M�MK>Ι��1nA+�ո�c0��Ih�f���!��Q3�3�;oEu��*G��(7ī��~~���X��G��&��(ȇEHD�;�GS�rMH$���8b˵�U�՛���4�
���.���K d�8���6�$���`,�����<L�f<��Hp�W����2j�7�_�K����4��xN�=8���1��I̚d��,�}Gw5�X�E�}��*��I2(������8��$�ȣp�P�&^���X	�f��`~	��PP��1�^ZV'k�,*�}��1����Y�>�ތ3�F��f�&)ǜ/�h�d\�̭CN��w]���K�����V����w����p[��c�*�5}{fm��:��75x��c��@&4q�`�����e�v�r�������Dpk���K��s�fZĢ��D��)����3�?�N��O�J�EE�[��������(򷑘Ȇ�+����g�@/L5h��i����\oM�`�����a ���������W5l`�9B�x$C�)]���FN]#�%F�X~�L���5N��lq<Р�fn��P\N��_�E2Sf?r?�?շ���<�W����T>I1pt�k�luSgz�z`C�j٬� Q> �"V�R��E$&�
���5�1��ܢ����c�����l���dU�D<�j|A%�2�����x����+E@�m��UqzBV���1���u����E*|ɳbC0�x��gu�9φ�ގj�h F[J��ۥq���>����<t�����K�p�;�C��}��;�-���%�
�k�Q=�ꦭ훨z�0(�Z���3��s+H��t���(=K��R-ժa��A�2������It�x�m Y�{�ߘ;��@ӟ�S.�S`��y���$cczL�eM7.�c^+��͂�ynƪ�i�v��Q'c%[|�}3�N.R�z�#��c�� �?�)x��-PtL]	u�d~m�W��K;��L��U'��P��蕕��I� �y88h٭��k��<i�G�Լ͎H�l�E���VWkS���Ɠ�ͿP�Oc9u?�~Bj���
c��f�z�=���;��a��0';`W���˵����["���ץ����\2�2�Q���;����BR�]���M\$�����Z��������p�°\;���Fϗ�wPט[R.	��Z㗗�Wop�Šq�#��� ��5����gGq�gj:�uʋ�§�M�א�%W[-�Y�98���� z�2{����?̵�
_a�2�T5��.V���Q�YE�}Y�m�GW��I"9a �%'�{2t�(��2���6��1��d~�fI$/����B�)G��7��l.�����
hjw
Yy��U/�N��+-�"n�n<I Z���QU8��x��#��_���`H	�+��&�^|X����m�_� ��$�8G��&���Y�ƾ 4�l����7B��)t�dh�YI�Wk4�2�da�93=�7�xk].md��-K�,�{�k]��h��[����94����o^	��T>x���_g=����ʗ�9u�\m��bԺ�]�7P/T5�`�T�(%q�
�ku�:]��7�Q��R��o�|�6U�i��o�dR~0:�=yn^Dz�Y�J��P���4�IY�yԬ�Y�/�z��D�ږ<��O-����J7�����,R������#��ZD����ő��ܡ��880Y�`�2��o�-�)��̬^Ǭ�i�#�֑�H�r>cDA�H��CV�뭄�x<���h�&i~���n�e�sB���g&�ML&1C�����6�� ����h�Q��8L�H��W�%�'�3�/E0�flm�����'��7M
f�����a�Z�2j���&|G������;��&cy&?D���v��y�g��g#&,��赍���1�D��
���r�s���0�H����jRl\\��_
^RO+|{>H���޻{��j{� r��ݦ9��";��p��l.�qyP���'�i��t�&љ������Ӄ��|��^��3�B(��p���@�o?��ٕ�rǾ]�����p'�"��S 0z0��E��ą�\r�6'.!9�ff"`ՠ�����'\�5��`��</h��5�L�6\���Y�!�4n��VԚx�D�B��j:$+��֝���t�_n��O��p�Ҳ�_T�YA��aBU
;��H��C1�7�E|�O2~�k4��v:Ӣ^�P�A���
�#�.L"��K�GX���]�GR��{~ sd���_���>�{��S9XU��[��������[N�p`ѐ�FW��͞���b
�$�
�빐{��dv���듁������15|�*!Y���jO�չ�T����"i:$
����;���ê��;Ni���6�)�GuT�3٧�}yw�&D�Ⱦ�پ����6q�%��iY�t�E:I�zTC�u㶘��C'��A�:�r�7�WL�]Eǖ��Wueo8o�dW>�_ �p�ج�Rx^��j��W�1t�d.f��/q����y�f���P�+E���;�����9��ί�b|m�k��+��!�5�4�+:���>"��n�G3�D��A�s����V��2���
����;Id�w^���1�Sk����$	�a��W�{(���c������߂�rA*��7�d�Ne7J&P.�/޵�)�.��KO��~|���"T# ���1�z��T�!��KG-%�S������|���9,*��M]m��!+�t�z�51�5�Y�;t�t��2"V8E���+�/3����㕅�K��'R�Ż��ǣ�'�[��X�FH�-�oY��L�㈼#�`���݈�r��:��ܖ��mx�RQ�e�r�H�J=l����̢<wyH�ܝ	E#����JFU�,�gK
Y�����K�����N I��N�z�\�E���C����]ZI؃��K�gy'�3�x���7"h[p�7c�µ��Kf�{�}1�����UGs~^'!����N8�t�AZ��T�t'>n��V�(��[��獹C����6�_����m����,��hI��.NQC���2�6��a�IyKH�M��/�{��|�d���Q!�ij�����e��e��жךֹZ���� ��Dnˑ�ƫ��pW�(�7��ڊ�1�M��x��h�)T�.C|���0W�&���9ҏwȌ�A�}��w��E+�TA.4��w}/�aK��ka�wVr���F���6�˩PzЍ���#I3��v����l&�LO\�G6���P��z��
�#Q���G�:ɨN�^�U$w�}O��_,öx]��/i��=���|S�T�{v5,�:\��E���:��Bb8X�n���u���b���IW��0W�q`͵
�j���XDǨŇX��i�?5E���J�-��J��B��$z��l/Jv��:��%���>����U�g��m �>�!�ej�`����k�II�ҥ���Q�$ٖ�h[�������(��au.���d��	N"F��(��Y�m���D��<Y�0�S�JP�i{����-��Z�W�^R�G%V�J��Px+��\"\������^S�J����5y|KixZn�G��lRXeOv�M�&Y�\���7.��.#�.Lm4[Nϭ�b��s���j2��>o��ҍ�i6��"�8[�_������#�eaɥޑ��4`o~��q�Rn*Ɠb�C�>Y�"�����߳�Y,��X^T:��	n>=&�_�;$q���G���D���%���-#%!� Kj�C>w#-l>^#�����~���֛�1nϹG$�A�����>��f��j�;1��P���r>W8�al��`E�;��mCm\{�Sײf�E�Q���K~�z�8ML����������Fe�\n�DU�܆�0��Z�j�z��d�АDF!g=R� ��Ht����F�.��lX��ü�����և�n*�M�
bX�� ��)�h���[�
���Ⱦ�Ǻ[��攫�5%�}�Np"�/����A
F��wPQ���=;A9n6�\�HDd���kk�?.��裄Y�[0U��=/��G��{������@q -G}�(?����I� %Ss��]|O��۬�Pw�ꮨ�5���i�|Ep�����z�\�ӱv�j1���l,䌟Q��3yDm��V��fh��<�?�R+A5s��ܑ����'FB���W�%���?G�(��׭���l/����w����:LBA�+��zO!X�a��4k��D��M#��Q |W���IF�A��9�NL}(cѹK5\����-�>b��/�}�Zܙ��5�@dS�d�����@��P��"n~�L��^	E��%�Ty��,���k�pײ�Uʘ�)�X_���T�hO?Թe0�W���P�i��}�$v����`n:�Q�
I���4"Z
��Vڏx~_옱��2�/�c#Ľ_�w��)��h�����([1�c�J�b�C+z�U��D�X̮���?c����~�SRGȰ�$TF*�n,���E.'��u�c��ug��79�ݎ�U���"\��Y6E�̍�V �n�gY�7�%AӳlM=�ԁ�_q��:�D�y��R�ヘ�PZ(t��.F���Eu<(�I�Oh���=��b�R��f��T�=M��3�>��j������[	���~�b��V�=Q�5��+X����Y�&~[���\\����x�".�����} wB5�0�͛�$mz%�<"�@g�a�w���MT�3�4����nl��)aV����Ȅ�RB��B�9�9��J���2��/X��
W�C�UN?��w�\ A#�^�#�2V�5��(n���$K��y�H�d+��:Q죎h!������wL.G�5��$^y͜(���������Ӆ_2�rx�&a'�a{N�����1I�Tb�X�v�����Z-�B���"*�ܐ�����`�����^R�Ԕ;?�r�P<6y���ɚ��[�ټw~���t��&m�z�sb;���ԯ� ��寀��ҏ�urI_���?�R<�<�V�b��� S$:���� �8���@���]1���Ú���ѻQM����l�r�����>B������#��d8�P%֖���Mڲ;.�1я�S��2N*����a,
��d�,ӄ+T��ߍ y2[��mg�Clԕ��߿�+���l�?'U�-0�O8��w�TR=�a�����x�?���t�U�Uw�Y.���E�k���	)�(1Ѹ�E�e#�K�,���+������+a.�Nޥ$2hP��аT�D�I���l�o'q�sf�w�r���A�����x�\c
Hg6�I&ƍ!�Gڼ�x�����=�s��h��Ĝ��x��uK��B�G=�Q-䯠��
M=ʥ�JG���3U�`�v.{�e�T�B9�h6�Z8B�[����	��݆�����	�tg�L�Y�M�¢�v�}s����8�!Q$�㝢-�	Dݧ(�ܱh�}.��BR#Y�TNL/C�>(��]D O(�l%��Fgj��݅e;x7��V��d�OЧZ/0�p���Yﴕ���7���ı����Vfм��xcI�xh�H�����.E��f7�3z2���h��|ʸ򯂝�=��n
v�gisJ+3�Rķ����k��[�����_)���'uPE@�Y�\X���@�\XA��E}�r�v��WGr����ğ�lf'Y�Zv����I�2�x��;�|�8QsB7�x0�Ҋ�ۄkb1�%����������O�Ȏ��6/`����8C�A�/�G�:�W���E��r!�@?1� +�����˞��_�C�g9�ϼ}qQ���͵v��&"œ�WC�Q&�G
/��$�T�Fm��\)T�_T�G�jL���R)۞��Zp��bB��^f`��+R�Y	�v���w�r��.h������{�!�W^�=T&O�����I�j�&`UÌ�8�g��ᤞ����|O��Vd�Z-�����.�)��Q���x4�H���H�������3�V��W�R��G�0����^+�����L�n>�d�M/:"��"<�?H���*쓔}�A+�Q�җ��CW�~���(*F>�Sn@+Uqc��W߭I	O��i�V���M(m��ּQ�=���@�_��]�%I�~t'�t<�A�6�5�z�x�lBA�5""�^�̞�罛�~KC}݀4f�p$k
�v:K���Qt��T�.'Øg�ڽ�.Z^i���4������d%��#��j���F��R�+~�����c0��R^��M�N�?n^��tD7�3��Q؋%��r�ys��E�Q��mI��}���|��w�)��>V�1�M/����̥xA�]^�4~ᘜMh:E�u��#�~=�i���W��Ӕ�>�V�<�UJ�����q����D����D\��ǛO�B�O��W��!��1�R-ME2C?��aqeA:p� ��br�7���J֬P/\���S���1�I#G��Ȫ��������z
��).y�
L��]�f�A�#��B�܊֥]��.�u�"�{.V�B��]L�҇͠�4tBE:�&�
��ق�>����� �^="�xR���0��.�h�����)&�H~o6�	�X���H��"ޫ��<�M��,�L���Ҏ�-�t?����t�s�H����q|sU��o�Ҫ�;PI<�Z�B��(��Q�.�`iB�Y9�p�X�Ǧv��Ž�T��܅|��H0�a���Hy]+\j󺫂�-�*�[-M�3;E)��t�UR}�1y�CL:9���,�:�6�d���	u�D�njGy��e+�X�.�9�X5ڕ�������z4����oy�p�ɀ1�u��u��)��I�[~{+���>��h������ts/U��Პ��@>�A;�<���	$�n��f�scq��p+J
�W/���>@W��G5h��e����Pj:���"I��L^��h�}�Ľ�ـ?��8�[0�!�9�� _��HM}��c��̆r�J	\Ҧ�`$�*��	j�N�$:���Z�H�UI�b0�����@��-��B�{����#'��8X�}X�2�D�Z9�b�X8N��-e�a[Ȕ�:����m2� A�heP3��ྔJ�e\�EzV�'��e"E��ĥ�+��w�^K�2g��-(��$y�\Y1�vch�v�ܾ�B<xU���緟zg��K⫪zR�u<���b�	� h+����,$�HD��0�NCQ�e����x�����3qZ��+!�����`��dG*�����X��֪p�,�֢<-ۍURY$`!���۸��P#�`/��q���.)���L��;R6	��/Y�`�۔	�X��ơ���]�v��F�2��(A�[���CeP�O��;pa0�� �~g$+t��
UJi���:uC�&=�`�JRŪ��0��+�'I7mW�{���������f��� �N��T�V�R
�U$V6���t����2`l�08��a%DH�&�(��?�6��C^l�[��;a`��$��N��Ov���]���1�|~�`ϡm� <Zj�פ.�&o���(v�:b����=�����sE'���ͬf�l�
�d��K��	IL�P��g5�^�駗�Ӎ<$�Å���{��x&:�ͫ�������vz�I�$�s� #<��|��6Nr�D\G$��&b�
��ʁ�y��n�8�yr�F[Տ���B7�f���}��
~ 7W�a"wתG��㬢�z��:���iį|�
6*C��E���|�cF��z���K=�'gk!+4L[h���e�^��e������Nc.�i�%Ya&z�pVOv���ex�\^`K`P����l9�4��>��F=��6��fd�#c��("��%�,���t1ê8�BK��Ŧ���$��X���iB<6&%�E���� ��ӭc���:�I���������2�i������O�e&�,��)�.�]Y6W�}`7꽁�� em{��;��xk�|R:k�S*W�����rk�3��M�Q[c>�с�ލnw�zBN�<O��Iu�f�7	tQ�A�m���@�臿��lh+��S��M��̃[���	�zh��+��3�4�n��af�C���i���@����ڡ�
�bi+��2����N!*!!K>�������B�K�|Vu� �F!WA�ߓ9A�eL��]ܵ�V�(��vf����_��J")�G�b��������U�wnH���	�M�_�?��:����@��X�kZo�"'N$�D�tCM�հ&�|���?��ث�[���wX�w�W�a>�96�[rfП��W-It^����l�۾�C���)|hl]*2[�8��[8�b�e�M𷯝�c��aZQ�Җ��H�?^4��u.��'�����z����)�ʘ�� z�#+��K
&6�;�>e���z�rd|��h�>5T�a1����g9�?��HN�jUr>ih��[N�\��Ђ��[qY�G�+�x�JM��<�r��-5b��c�[4��\�������(�}�v{S֪�Dsন���-1�#:L��lg(zD~f 5Q��Q_�E�]���\��#	�k�T49!8wk�n$�.��2��Ч��-��}V�m�.��֞����L�89������:3�w�rr��ok�8��4t�{�KF�d� +�^\�-�`ǭ����ͼK���Jk���0bq�5��-gG*'��;y�)�*U�M8�=�',;�h�ϥ�7��t��1(����-����	��3ӕVx���`�������r����v��CJB��l���߼m�A�7#Zɤu�Å��t�}jOԻ�lO/5�F���uh����s(�ښ
�&�`lw�I�0�a^�'�?�Yº�!>!�9���o"u�4��II���l�����a�o�fY-0M�����3T5�H�k� ����ǌ��m&��ͥ>�o	~a���\�A�|+��[{�kő6�/�-6�qF_�>r�'$�_J�E�-������y���e�l�Ѡ�ΤD�(O�߶��Pc�"�`=���JH�M���Ŵ�LС�QbP��X�#'�~�?��Pp�ǝ�u���J��O�%L(�E�V�S#���7�KPG=/+�w�Lvc'�?� ���
���X��n�'���W�˽��3~����7��� d26��'�M>�܂.��*.(��ᓛ���\�e:c!p��457E`�1Q�SM
� ��h}�ӆ��;��\�t�2�o��n7�g�(r#i���L��p%y�`��0e�u��^�;�@`�_}�*�pq�IA�ʹq�*� ϒ�pz���x&�X}���`�Q9��	z߫{F���#�+֟[!��؅5y�?��Wk���M}��f�{W��\���'�k���\n�q�AN6�̭����2Wmr���l�;�b���#RZ�8.����= �c?y�N��SI��^ZV�MJR�[�	vbt�!����)Y����X�����̻x���w�ƄoE�m���RU�m�ż��"
b���D�(#ѐL�BzGI4���fn��W��x�gu�s��E5n�Ć��K�^>�܊����`��+��n�� �UUW��C�<ҐN����Q�H yt���N*O���,d^~�HZkA�az���-��Z�-�2+Α\o�q��:WT�^�sV�C*	��)�53>��Yѕ���]����t�5�T˲d��מЇ�?&a`��U��í7�����0[��ݮ�R-�;������.ҾݙV�x;M/���`q��2�V�B(��>%M��4N�qHf�4�is��Ā�l�����B�PO���_�c`m�GU��,"��$�
Wߟ���y=�C�%d�\�=���>i�)!�3ry[�����C�fğ��-�{_�7FO{�`��=���x��v�����`��=�_8���>`E�����w�c	,��E!�'���匷VJ�����މ�k�[6R6����I����_[����Õυ��*320�Ln%�\�B�w���pi?��.�Aޥ���*��*��ş�G7M��>�����O�m�|��Ϣ����C6#Ϯk@b�2_�(N�H4�(uf��,���OJ5T���B)�I�}_�[nҦ����J�g��M�U7�?Of�8���j��!�̇��t_mߕ���w��^H)'�z��W�<i�I5�z�F,������_ݎ�p�tk��"��� "����Fpf����Tþ�}�ϐ�@2�{)so��vd*���
�+��#zZ����?b�@�y)0L��0�QF�'�$O���ۉLX�M�A��*�(�ƥ��V�֎%�ȷS��L�`�jLu�[�M
���B�JoA�D��,��F��m[*�#�n�J��i׸�	^�>��%��Wo��oz� "�M����!�<���{L���Q�����il�	��q��4�`�z,��Q�[�4�����fŠA�O;9f�=Jyet^�^c�N�%�;a$-���B���JBY�b�ufU�xфn1���M��FC�|%�o�8�f]]�)4��T��9�F��t�\;��'�t��50I}~@�������Q�Y��lx,H����+�u�wR���)�vzJ�˙�n�[H���]S�|{ @`5ț�ߒ�r�8����ܫ�c������, ��pp��쐐���sR�p��j��LA{�J����6n0g�ÖCΙ�S:}�R���S��KòS�" @p2����;�ɳ�y�_��4�b}�1�f�\�Rt�1�?��W*�	&�)LJ��{|d�@b�T�4% �BX�4�� �o&�n�v��.�/.�x^���jK������D��\����Im�7GCR�|��(7��8$)� 鲆㇐�:��u�D�%#T#tr#�{�ԇ�<��	�8�j�4ь� ��R�PJ�'������}�w!L��x-Ҍ������Y`�irI�9��U����]atx�B�? �W�^f�}�$FF�<]n�}� �a�b��i��}ؑ|�Z�$S(X.�vn��������+"1�W^��"��U�s]���^��6G9�>��M൴� Pp𛟕\*%�Qm=c�i
0����7�{�l�寈�z���!F�_>D\@TZm) �GIwYEG�2�>X�^�+~�|�����ޖ'����U�ܩ#v�}��P��oٜ]�R���É�B���ǽ:�J�Fv���Ի?�2���!է3;�!K��gmXbuT��7IԊ�5�m(�JB�6�G�2����ڼꃀ*$����<g	o0���q<��V��j�C�}=s�+@�}-��u]ֱ_�q����4(��s�Ĝj��T�]�0���8�8����I�y���ԽK�J��h��-��>/C	F��r� ��y��I(�P!OT��� ��ۉO����W�V_������%ܪyB�\�|[��_HX�}�Z�����I��S,"��0��Q�C��cF���� 8�3X-�3c��J�a�_!D��NÃ���*v=�9[�YM�����gap�w�{$��J���N��4��mF�;#�`ȂbO}��L�
W�Q\�m��ȿ�b��s�h���ʅ�􀱗��kJ#�鲐��O���Qѱ��v���Y�	Jw �>F[�x�X���Qw�����ئ�P�=XXo{�����%8�<�t�t�8H=���!1�4*�A�c�r�
��-2��Q(;)tAle��6����VoE+w�Ȣ�q������h�7�� [8�\ޒ�We҄�Z�pѴ�]�ݷ�n��@ҚĿ���.~.+	����_�
��n�^���9��~������LbT�D���̂3���&yȅ�N�?��_<{�[p�����r|A��Է?�?lm'M;ōt�?�r�P��'Қ��5������t�Di�h��̶���YD�sBw��Yl�K�{fM�&�Ӯ�fGՐ�U{����K��@�D��㫃*'i�h+��#?Wڲ�W��<�TJ'/s�@��G�UJǎ���;�r=[y�	��$�΃��FV�����Z}��5��ѵ�Ǯ�(�>�-��t_���-���d��CQV��6��5�"�~6o��b+QR�k��.$�`υ+x۵ۺp ����PX��v,���e�]d���Gqt�&�90�N���$^��,����>�i�;9Sz�6֣w/���Or�bw�0�@��:e̺�j���:C.���9s��z�E^����*��c)�FxA*��j���(�h-]��3�4�|\��h�j����4bm��H���ب	�����󣈸t�s{�����!���u��m�c�/�g�hpnA��u�Ѱ�"��ad���G2�l��"}��'6Y�
�uE'�p�y'F��^aam���xt�|%�&x=�F�5:�R�������$tu|��;zcԭ�ݙ͚�v��&x"0+��%�FXFE���L�C|��U
�<� Z���v�ُ��2�8��J��a���,�A�ӱ�������Lx�#�	����S����?�Fsj�sQ�	�#����R�ć#!.I9&dX� G4/��@?QHڛ�,D<���Sd���:n�K��L�$q(���j*�V�j�$�G�΀�����i"	��$`u��e���.J��(�+��]i�3�У��,>E}�C^�[��+M��6������4>�8�M�m�L�
�ף>w�J+���bb;
K�@w�R|'�.��C0�U�K���q�0(C1�������k�?*�#��`�JU%��Xo�Xc���L��ߥ-|��H�>��>a^��|bjj�
�ȭ��x�_������@���k�/��������g�����<�jk���Q��7%��>�S�S�o��A58�v�!L�Mߜ{�h��h,��r��S��?���������q����jc�]�F��y�*l|���(��������O��"�HAW@1xSv{����#���)���j7�� �Nf��)�/���=���X�N
7����̞�vAB�bp��D��;?T��5��d΀�{�j����jM҃Ј�#�g>i�k��sk��~�.cQ^�m��㓠�n$�m����n�
�/�ȫ��?c)Ra9Y�w�!�wn��5`l�w	�fW����{s�x��mRǗ���͙���#��;:gHW?GJD��3T�S�JD�"����,�ވ�Ʊ�g	��wK��ˉ��n�k����=�����F?�L��h�el�^'�qأ�e�՛�n��g�ǒuB�[6�[$��-��_(S���]?��2�PF<��-s���|�����S�̊�D��b1B��R����>�Ɂg��0�I�bw��{^�N���l��V��:mX҄�;c��C��v$u��O�5a艛͐Ҹ�L��t���Tm��(���Eb�$�$�@-�l�}(���zW�Ċo~�ϊ� R�O��gi!lj.H���(fψH_����?k��㢎zpR��=˃�ג��s����|O��#��l[e�
Q`a����|rUs���jf>��Q�My���vE��8�_0�^�^��FLQ�D��}��o1}C�cW��0,�����
�bb�7=���}�7O��)�h̪��.RU���&?��a$sz=S�B#�j��qj/�,��W����Y$d�qi�"/3�Q�#�<fD��a���b0L^Ɂ�,��pC�s0��x�hݽ=��hŎ���[� a=䟋��B�NxmޏZ���]���������� \@�Ԧy���n6󪃙�Fxd��B�6�jB<�6��ҹ�ǐ�0&^>ܭ���Π6/��M�k���4�h
� ������8��|�q�*W��}K�Ճ�ަ��2���0��ww�~r��/X8~�B�/�^.��~�z,��J�H����hwzS�+Qr"O_�X��cR~@y0ங�,����v�.7��c�*��hq(��a��e�rh�45��h����#�1��T�(m��0Y�N4{<�ࣺ�䎂d�sY�#���������׆yB�{�|.�-��ʫz��!x��O�C�}��:�>�� ��7{"b�M�5�m�o!)�B�"PϨx: ��J�Źih�m�{@ˌ�dbkk�4lAnZ��6'�EPdP��3����bCR�E�g��!�v�-V����(EyG�H�5�!�JK�K�������w>�:N(��pN�7d;A��ޏ���J43h��b,p�t��b³��R�R+�������������ZcZ���#5f��=J"�m�ox�%��A��qT%{��;rN�@)���9�)�F��X :�� K�V�0I���l>CD��^�B
�Qߙ4{ƺ`];pB��+$B�w���Aq�FV�K�[~T�#��<�T�|,���|u�kѝ{� Ԓ��,��쭹��?/F����PK��"e `
�{��&�Uh�:��o�e��3X���L�3<h{�n�P�tc�8���#3�|ng�s��_��e��6�[�n1�`������f�9f�J�r"\��6+<g�b&��b�W�;�%�7�ҡ׭��O Di�Au�ʜߨr'��pq?d�|��U뉔��j�l���������Y��cˡ�_�L���Ar᪩'��k~�x�	z�*�=U�hy�4������;�jJňO�q�e^D�XX���[��]3�lCbbIf��j$�[den�~��hz��ߐV��/�m����/����K|D�C߸?�W�M'U���Ft�žT�L��Dkc��	H)w��A�3�gf�&��	E�!��K��)��$������ʎ��y���'�Ϣ{+�j��"Gh�dl��j�n~J��F�ƲTE�$�
�����fk8Gݢئ:^(\��s���L���H�xV����u�Kԃ�R{z�Ѹ�o�#�ĉ&	��9�1��x��P����`��� L�I����(��$��*�ݽ��ȍ���I�E��������	Z��۶+�c�
�p����=�=h!ٯڕ�ES�!�6Hcs�:oLi�"����� 	����M�W���Th�\i�	6.�s���h�.�[x^�����^m�eW$_ݐ������ �is�$�)�m_���D}���*��yT��W���]u%Z���O�d�)6U��ra��Ȑ���:�m�BW��xW��0 �����(������f�OmA��w�5���I���+��tc����-����Đ��wSf�T�]�{�<p/�ʿ�F'�Ya�~�6Q-�8:�@�����\�@�V~����ۜ�=X��;6�)�TuH�!�rƈ�ж[�Gq���u"�Ƴd`H���q'+��̆.����3���1EӲ�̗���1+��B�E�4�`�(������Y��V���L��r�Pg5�BVH���&��zFձ7�צ���������	�P�|��G₨X�	�)Jʽo&�cV�2�P�(YdO�������)��dJ:i���kќi�j�<��!�����@��%I��;t�=ROԄH.�$+B�`��1�g6��DAf��g^�H�����\�T������9;�?,%�U��Z�X�,.��"�q�S�%0���%o:K�U�Jt�3t+���� �U̴+�H$y9
�����\�ۿ�u�@��Am^e�WCm�����9�z�XW�_��l'�) -����Ȟ�qI�X��-��C6B�M�)CS@_��
���G��v�d
���)h��ͽ��I �q��f��aN�f���4�������xh��j|e��t��qlQ���Ff��l�ܭ��:�\�N����f�&3�?Ck��5ZR�bu_B�(�k1"5~��&�\���hi����n���{:A�%��>�h����௖PRF��g��˴�9��N�c��\_YC��R_Y����Lqǰ��1;�Z�4sP|O6j�ۡ���r��Ӿ��Q��t�*�[�-F��inPF�a�r}�����_��z-�Y�3�Զ�ōfgW_�y��3��[O�����ȌO�m���mlC8��x��2hwl�&�y�H�TL3���8o��w���R�[~�.U"��\��������.dڦrXe+ �D���_\l5=}i+����]j���~m$AK��t$Ȩl��'��*�R;��Up(�p�[خ��q��0�{����@�F�L���͖�ۧ�\:)�&���Qz�� j��M�����j$p8<5<\#��,��X| �Nb�.,�A3������ۄT��e�1(I�h�M�`�Z�ΩU�����'�g�'z�}��yA�;~������M u�-:Mi$��{�q:��à�����S����_b#�h�?�����d�	�����!/���UM��yQ؂N-# j�*�_ӛ����˷gҢP�M�����0뽁��יx2l���W,�#�Qz^��IJ�E׶J���r��Rs2�&�G�b�&��D7|�y������q�)���EV�0+�/`��Jb�[ �Ru���`::3<���0�I��U���*����<J�b�ݗ�糧��S�)��}u���/�ࣽ��1�>d�H�|�k�������|η���<;NerNkS�?3�^h�y�y�)d��@�����I��N�}������w��?u"`�ܞD\w��s���,�@����r�`�|7>��6�sF_d;|$��[�w��i�u��t9�>f��?K������k�;۵@@-ɽT�nh,T��Ǿ��뭸<	WCWY��,q��O����QQ�0h���ҵ=S�o�x;�s�Q��@9�W�ĺuB{��YҎرi{4�A�᮴�v¼}U�[�ɦ�1�4k$���#�J�j��}(�Md1 ���E��G\@�r�DI�Q|ql'eK['��O_�Xl�Y�u ̔�â��r����g��Ϋd��ѧ���@"*ڵL�{�k��Eϣͯ�SX�
DyىR/>;��.Y��kzR!j����}�µhK��>��
~��x�?�V�p`�\�jV3��*��r/.������AQ4|j�2��� �������G�wڔ^�)4��UZ;�'�:YG>�O�9e��-G��\OH#�x�mNK��<I�=�F�?��E�U5"<�LV���%��{Е�]��r��s�,jKU�//p*�H>qS�4��wS���K�$�Ƒ�=���g��~�\�� �.9"���({E2�W��*���q7�听�;u�̞\��Kc��|��_��8�HMk�q8?�!{#�9}�Q&	ΙR/�8H^�!R�G��<Y�+Yg6WE��yI�I�@�ŲXnb9*�4��Y�:
�j[kFE��E���������0`eL��^}����@�g�/2�!�S�(�B�]�CI��0ݯ��$��R�B��:,Q��r�08�Q��&^�)ހ���!\ Kc���?5��k�<�̤�;Z)��'K�e����l8��G����\s�,Q��E��#���b�m�ZX������/�eM�Dr$��2"��K.u�~!c�-�;�oVyK������g��P�"f 8�/)xD-1GY���͒���a�/N%BH*.�^Q{<PE9Tn�{<P��&!�{@���5�!��Pw�c�
�:{|�� d���FC̽��ɘ%D�S��F���5Zl.� �"Jf[�����#m����F�`5�%s��ѣ��Z�����7��F���^�g7�3�|�os�z&���f�7Ė�<ұ
��V��}�$�yB�BwX���L�rDL��3�n�2c��:<���m�,F����|�  _��&ܡ��]�^�kUS$�_��<�3i��rg�g�z�>�> D��U�jt�c���3#U~@ZKE\LI�n�X��~��t��I�.�d8.M�y.(��t��@k�{}XY� Q��b���Xp�v��U�J�DGY%غᆿ)��T!�Q?�������Ʊl���uF��[��a9eA�fǺ���&�u�X��/Ϛ�]?�ZB.�!#|X������)N^��Wk�)U��e���HI�B{�X�0�,�����p��r"����{�T-�v�[
��ȇ��;�=�E�nO�����6p���om�f"�IE	i�" aiz������oݙQpҕ�L���}&%̈́�j��+����&[���H�*#4�d䙝EF�sg��тO�*D������Mdل?���N�bL�^X5��CD���=9��}��I����|��%�T�$ �G�!��H�����O��<���֍�U_�0[��nU�]i���AR�)h�M��"@7d4�a�Q]�Wəm�V� aN��m��'�&\�e8.ٱ��G	�����V�j�i�N�o�=��d��>q�l���S����'��5":+��JzLRn
}�3�W�_'�X�)�Ƌ�Z��K���	k�'4�|�HX�kE�5:���Z(���Mc�A�
F�m�y��>��WW�v�o��,Z��}ϑ{�tj�(����	q�,��i�
iT����b���6=��4b��槶�ry���D�l'R/G�E��$���������p�֏x�`�sD�
*z~��i�/U��u���4N�Lf���fP<�]��2�z$����:E���ٟ�Ql(C�A�c������[�h�tZ�l�+a��ƭLo�3�
�G��Ҭ��\#���W�k�r��+��W�h1+jV�%v>p���[���	O�D�\VD��������3ڤ�Z~�"͸<��Mg�y���^-��D�Xo���g/�5�\>�7��Ϩgu-eXQ����*)\qư[������+$<7~�4T�b�Q^PNz:]<��`����s���G�ʠ��"k�l�
4a�f��3���'�_'�{�(�/|�@y1x�;:�K���9W ][m�X�s���!�Tvsr�+P΋p0"�j�t�+���e�͙�S+L�(N)l<+/`lIM_�d7�ː�Z���&��B�&lk�"��2�`�m�\�6�v+�P��i�v�v����;B�nD�ݧs�2v��}kD.���1�����|L�l��̰3�rE�Kfbq��)Q����؆�#�o�����kq�!ŗW�P�2smk�����=}��T�44&�3g�a,��TtT7aj����u8�����O��6�[�S���`��WB���������>�V���/����;X��;�ɉ����w���]�0�d�0���c�~%�S���R�K[������Fk��埳��F���ff��`�U�!�*�'!.敨��\�$G�ñ��`d9]er�m�$v�� ;�2r�k��"�3�~���nl���{�tm���,C�,�ʂ�[�G��+I�gV�hd�$}ן�Pw~i{�m���n'�*��`Xx��r��$j���6dY�=(C��b��I+A��0�8�$B���V�f��Fv��k��Y����!��G�བྷ���zF�E[�,�K9	{"w|p����7yK�W��Ƌb�:�0{���/nr���x|t�?��ZSa��s����a!_�J%���C���4D`#N����;���?C����Vf�:�W�(I�[��=�W��O�rd��þ�%�.�H��G�E �[����8x�͔<������Y6��!7ͅ�j�l�"��#��jX3/I�nᵁ���*��{z�^	�O1�6!>���aQ;�t3FY�g�+#[L�4^���jpF���Qv�I�B:��0�@��:c�{-�J�bw�~�bO�|ǉ�4�~��)Ӎ� {��4����$� �|_�k���F���!�5K����J�6[�b���2�`a���Y�L�Qg��=��K9p�bf�?m�&��i�'8AÂ ��prEΉ���Xa5�r����@�-������z&����]����n���| 9T���v����\J�����)DeiLPy��R?�mz��N�/���QLFw��������L]aωdZ'7z��&���){�|�|�o�?Kv����P"�I �����Nl�`<���-z��|��G��&o;��b���\�&F�G���b�)�]}	�Fq-Y, y6N(�0� Y��������S���˗R�v�
(�����Cն�n����L�{
�
��e"����f~:���
B�l�x����*��Z�w|����=T���pD���?�bi�}� ~!�*���CAAg��p}�^n�@ڨ)�'?�E�����n�#X���j�t4��-B
=%=_�t��B@k"�t&���6�g���u�D��=��Ƽ~���j�r��mbSxŵ��&F�]��j�K�t�3�Ўݭg��jv˼��w0���\@�uӾ�'�b�ޒ�Wh����t6�V�	�B��枠7�W��!���2�=c0n�s_[��G4�.t��P��?B�FI�YtߜL�>5�=���r�Ƃ�-�L���$��o�)vӟ
'�Xպ�S^\��+�^:�DхJ�-����?��A*"/�ᲬP���I�$p�tW�k�R��U��!F����-�U�I�)sЏ�9����8k;����}���i-wƝ�+�W����t�M��˃�f$��\q<f�7�j�r�^�V���%�jT�ßS����k�f�s��FG,I=�X{ב�|�� cB��XI;�QH�=w6�� �B^�WR�w�ʸ j�"�dZ/�7���q��>p�AV���w���+�9��;ag1_ß�ʥ3('±��O�RÌ?'A��P���1�څfx4�G淛��p��ϥ��Ju��[�;d�N��0�4nԬ�;n�ƕDЦK�з ���j���	I�1Oqu�؀���i 2�fXn�e���N����b#�^����=��*�a�t�{���6&��=Z��F.�v�l�M�o����.���Y`��@6f"UR:Q�~�E���Zd��f:_�"����ğ]���aM���'I����O&>�6��7.W^�;�7�ʭn����<�#zM���s}8��PN��t�U<T��~�^�sٲr�cjR����J܂C��7<l�S�!^���(8�>{l��$��ٺ���j�M����>���x򥘪v���F�#��.iJ���;;׬Z���ZN2���,(f��T"�Ǻ��D�$+y�wm	{�4�HD<�WZ��ϿCﮯ��^J"�|��}[���R[�'���O��;�	|���.�%���	��W�2�Z�ʧ�F�[�;F�n��|1�&�ok<a���N.�¶��:%�G�_	ѴHi�wrIY��u�`ݯ�#(ޅ�:��T��{�w҈�Zj�-$�'NK�9��3�֬J�m�ض�ҳD��F/���~�~&�d�1-�Y��	5��8 /��5�`9Ȇ�=��
�9(r����c7�v��Ź�#}�,G�hG �p��|�{��i�}�*zOO|��S��ό��k�B�	.w[����/M�e�pf��+�R� �40�\���Y�yv^�n�Ue0 U�Z&�dp��L���@}�����5R,��;!����/B�/u���x[sL�z�
Y�&2��s�oH�nc|g���h2r/٢�k:�p��x�
Ԁ�:�p��_���P�}���C]�7��6_s��^� �xv/9�+�Qf�o�4	P�fb�X�ҁ�K$�HlKH���}�y��'}��_��g�$��!m�)��S�Ht����5\bzv��2�ќ� ���n���1Bv!��h2Ϧ�̩�|<Pu`G�\�y<�mAf-s�B�v4B���,�R�!�F�8���o��kC/���3�M�vj��x��	~�
�d��q*���n{�K�ۦNj�&h�k��(ħ�VQb��죛�T����ϥ��h���� ���b�� ?�[zM�Q[G�VO�z���/-l�E��[y��!X%"}1B�����>%n�P��#��%����V�\�RIά5��e=[ifM���x�=�2N�O$�t����;7�(�-��|M�ӣo�$�ʑ=/!�%�j��Lt�h��`_$��Q���~���٠Jj)ΫYX�#�):m����,����ުsMn��Ho���CZ��q��'2��A������HR��t��J���U��-ԯ�a�<��"�c�ϸ`1ͺғ�9�@�.
mr�Ju��qq��@�y���6u���鏥E���ĝԑU���i̅2.9N��VSa�XU�`�[')��\� ��3t���ķΛ�4 O�g������YP�b��s	#
{/����ߕ�|=����q�p�B@q����ү�؇�������7��ΰ��:��Un^���k��������=E���_�,��C�d��`Е�Y0��͟Mu��3��:��q�Ɓ�MH�u��������g�S+:��� (�e�쥛(�7�Y�d��GV���ܳG}���ީm�^���\�)�#V�8�����΍���P!�z]�F��o�`t�x}Aeʇ��y@��h��FQ
��MI��	�I���'�ʜa������z���h���K���"8���t������sc��8��J�:��G�m�+�}Q��<�2.:5-g�<����
�t� z��21(_�Y]��	'�WL���0���K��MO�-!�'�\>���"�����h�^I��,!w��&c��L����Rz�y�j�t� F�܋��e�B��_9(1��W���w1&�L�q�=x����Z!2���W�=7��T�Gƕ��z�<jv�K�A��:1���Ey�]��z{QzX����)��*he����`�M��
J���,��4�l2�FAAW�±>�Km�yD��Z��u����iQ�^9�V�
rC耼�\�Z2�L�@��c�W@�w�>��g�{m���"��������2ڹ�����	'*�����3���~B����}A��OZz��Pb�\���
���U��$Sޮ�$�b��b��^��ER����@���n��d&� (w.�P����*�⒎�Բ��f ���7�Q$M�"��� M�@NȮ� ɒV��#��fyS'����dV��ki߮�L}��U��&L��8��̚&��V�E	��&9c:\��=׫�G��j˝�*	 W�[<����.�o��c{
�2��lIsG����ޚ�F�1�HKΡ`�ܯrM���?'�]�����~�_İZYȶo7�
�w���#i�=SH�+�6|)�e���A��2�*�ه�^P��.�KF�?,�/�5�vx��M������Q&��f��5_0O��+}R2=Y�JP���z�J����.�M�������1�K�3�������Q�ɽ?"� ��`��s����]�Gb�Z�u�^�@B�*��?6 RCFesr��� ��";Ey�C{Y%n�E����deR
3`�B��T��2�.媼�9�5��e����R��a�4T#l����Q�=EjC��R�B�l�|��
�13D_V��yE��V?��!��v���]�_��O�j���  N�����zJw���uq$���H��"�1:4��	�k�i!�bf�D��Dʴ�)%�&9W~U����=Q��C�ʈ�
�M��$Z���,P����W�~�������(�>!0xt	s��OGC��h�E��C�#O4�H{@X��F��JE�hF�#U���-�h~b�s��/�,5���64�Při�[�����9m�H���T��L(%S]`l>JR�_�g�������W]����]</~	[~C�������7dX����U${U(jT���խL#���E2s���7�)���pN�D���ӿs������f�i�yL��C�^��1��\V�*�0�ث`H̫�o������&y� �m�}���Zs���D61nw=fP	�H�S�Ȣ�,n�5�qK�.�Ɯ�<f�����U��g�gsl�b
�E�/�Y퓅.I�a1f�x����W��N��ҳ��p*L��O#ǟ�J��&>?��C:�;��0�{�9����)��K���D
CA����A5��ʼ�b�^�ۡ/����Ҹ�{R7	�H1��o�'h�gփ�
��,��<�Q�[l�N�.��X �UK8L�3N�����a98Ħ!(%|Q�)�aфc#F��#ʘ�Y�$���Ov咐��2t���<˼���;'�3��7_�am�		�P��@М���36�X����Hȡ �2I���q>Ͷw�~;���@�u�hs�.����a�3��� �����;U����]��[T
 a@K/?�ҳ�&�Y�<K�=[���Jiw�7
ސ�Zx�"Uz���ۙ��]�|!I�<\<#�����0���P�ۣ!���#띦���V��b۽:���>���P1�{���(�s����t���!�~�@�oM���7�TϘ�N2�+/�6��V�? ]H��:�EC>Ԑ���(a�T��x���
߬c>�T��e~����\���`�(`��6WE��;�z�i�eA���B�@Η�+���r:�!������D�#"�8�T]�~�o�;K��S�E�l�P�K�Sg���8`�cʳ!�M�/�1�� �	�Ηd���/ɖ���'�~��0�����0�,'���j�S�� <Lzכ���ؿ��G����$����a�~����H}&���_`k���t^��r�o3�ٔD~7WY�6�=��W@��^�j�E����?x�R��Ƚ��� ����g?��㊤`���:0hKN�7c60�e�W~�6�K�/����6KSJh�բj1���;�M�%��&+S��˗�܏���[���K��.jF��F����#�w����)��{(�N�h.�!v�&�&�R�0�	����$��K��7v�Ψsp�S��}�%�)1�vPF$��Řv\϶vi�A�j	�<i��d��3	��pf��j����'m�_ni��2�KUg*v2";�<~�ǅ��|���JE�p����YK�W�<t���� Fs��j2H�sj��� r����]Qmj?��0ae�"��rCS_V���8*/`p���gd�f5|�������[> ��0���%�ku��:u0?w-�Oq�BNZ�Ƌ��9UB���i0�QJ@�{j��2�>2�Pb �<�����k�Ҙ�>�����F�i�a�bj�i�b]2��Guy	o�4��?\�_�?��x[#�U�}Y�w��3�l����;$�ME4�.P��
�0KE|4=Tlq{���J|e	T�\|e,\,s��N��7Sx��[��=,2l#���$���v�����G�R��5T��Y%{}��q�[y��ȯ�;�IP^C��~�
YWk����G�eG�Te�ac���<��4=~�~�[9����ѝ3SA��{ M/i��A�ҟS�6�S%��5�^I��(x�������:ߘ�{��>�PEUv塀��]3�xB��N��`�L�\Z�%����._C$ٗl!iNv5���=��pdw�������62[r`�TPr�J��u�ty�+;��&yY!��0�c�{'(��Bko�D�3�ay1����驫����إ�և�8�&��E�Rc�P3�1�
҃��s�E�F�z���A̖+��0yG~]�P�v#�6-	-�Fx�O{�7z'J�Q[qk~�W �� $�G%[�D���l$��x����6I�yh Qh���Ș�����a8��_���=�l� �H��<�-~���4]WF��%�t�i'ȖI��f�x�mc�|> ���\����YF��7}�]�̬S�T_��;h�1����o:��3v�($S���g�����Xe�|!��'Es�"'V�$5&�s��&7��G!U�[�Fgz&��D53�Ѐ´1𤅰�4�*�3RuK�׮{F��魆���Z疛A6��vǭq�Q�j3ּ�4��}(،�+��p^$!�BhN,�(�u�*�"�=�����!b��`_x��R�&�ح[��#r��[c�>}�B}-c�H�KWγ�ӯ��?��e�{v�J�e�W�_i"������y�K�y9��3G�'�KdG�I.�B:�UN��ߛ�X�;U3��*ݛg�vd|ܘ��=B��E�n)�F��{��l|�r���QsX�|���2�"�ܣuk��R�q#�H6�ːt:�,��]�B��|3SQ4s5�?H5x�#��c���g3Ŷb˖ݢ�@���x��G�HVY�oo�����`Έ��y��f�%'�W�d�T)E|�K��3R�Ә �-h���@e�侚�n��X�2��Z���o*dba~0y����ꍨth:�S�q�OjV�[)V�$�'O\�m_�R+��w��	�ڭ�de�4�m��S\�O#�¯��ƸS2�E�$�S�9��TyD%L���tgV�Y�o!�|���t�ZXM��Ij�ݞ��3���U"�7��������۶nx=���V�3��'mx�����I�_�0V�`�S%u�=ҳf��nN�V�@L���"G	v?�غ�ط��n
ډ(F�]��?@�]�7��y�i
Y����bB�t�c�ȳ��/P��Ѡ3J�ؑz��n�ʻ͇dX7\�9�:\^�P/���~a����*E���n� �g�4/V����h��Ś��n��*H4�zO��.��Ά.�lLt�>�U��]�>ϝ]j���B{R�2۸�/���ƳF��S�K�����o�쨬H����J��|�_�	r������jicY���U�{���)��n�C6�C��zU�7D!�B����w$}�4SYCR�X��\�"�Rp@1���# t� ��5�/ M]kݘ"w~=���@PFY��%vZ��������m��N��s3<՘qSks1�w�������m�|2��c$ڕ��VAn{n	��s�R*�L��OS�_A9��R��c��7��f��]��7���[jbY������kԹe����7DHVb�eY�f����#�C��j���� ��A�=K���5�d���{<8��D򒉩�h�(��)�m]�IC��zbO��QQ� �Kq]\33�x�O��$s�*2���!��M�:�=Q�)�N��)ff�'����ByX�h��u�{�J3�ސ��7���P�(��"��t�(󊥯ĠQ@ަ�Wi��>��S1�Np�x��W9�G��\��w_׏:L�t�q3���|SWJ(�j� c��k�� ��c�������I��WĪL-"7-�@�'���%���ϭ��2����-\�ʬ�7����|��T�q!cNQ&�k�>�(�* �*�6au�g�-#R���-Z��b1螙 ~�~#�ƣxn[Ρy�>;������bBQ����#{�����/=�4��$�ZB���J
Y:4�Co4���.R���|� �s��zk4�� �vr=���KcY�'�q3)��X_��xu��@��D+��2��ζ`)'�@j����F��ʫ�66x ��7*�N*^�^p�EJ�'����*M>��8��.è:ғ���GNËc���(�nf���Y!�Y��3��N6�i	)���+Ўq�����<.���V����N��:h�����n �'��i-4���~�b�0��.�]�C��)n��q�߇����+���/ '�7���K�����ە��"��mL��~Pp&Yi�C��va$���d�m�A���}�l�uZ_�чΚ�O��٥��rʙlPmU[���4�e����;fC�<;ץ��"����̀�m�7M+
(븓�7�;*���9�x�д��س�Ek`�."d��lL�����U�ػ?�cRu�*��o��1�W�W`�v
������ˮ��r�����CDF��ӟ�8��lmU��q��|>Pq��L���
�F�q�����Z�eO��Q�एu���#AQa�؀�{&�[�i{CU��B�Ѻ��2!&p@��ғIR�����?AȊ��Q-��B��n�ٯ�!�z�:7��֠���ޥ�#��8���a!:������X�&f�*^X��#�m5S���R���_���GK�t���7�o7���<�t��EF�\/�݃��S�$Ȭr��ԟ��-Z���W�`+��1�Xd�a\2�'��.G��Y>l�ڏ�6�>�ge�fKy��)�՚��"�&R�0bE��벪��Mz��Z��v]`��x��(Sy��i6����G���mU*H%<2������WW�D��C��wcػ~������)&�����I���y�*���C�T��y�3��?7�k�4`��m�`º�l1��Ҟi��Yxd�8�4T�g9���!OvےF�k���p{�a�V�mu��͔֚1.���1�}^�B:������r���JJ;Ӆ<u�ܸ��<A�}@'"�=�$��(4��gA�;em˹�Pi� �7,8����SMЈy�*�f�`϶,^&��ju���`�Rd�b/�*nxh�i�����F��u��<��w�G,��S�f��M7O��>�˽b��s�S"raL�vb�~�SN�pz��MƹO�\>33	Q��V���wx�#���'�O,\��9?@��2�A�R���ݖ�|�R����:��Nbei[6��MocoN�꯷*W�M� _axZ,&���bi�>	hwf8�*�}T|s�ۈF��).�<��{.��ꎥ��+ -vn)Q�S�����W�;�l@��݈�٠k�	D9��P��+�A�����X�D��^�1\?w�f��gۭ��G�cTy�>V~up-��*�t{���:�_eXE�����q��/��a�ͫ鷛�����4�^��	���:k�t,���n��10��,԰�m�a
,��?qɳˋ��"���.�p�E�XWS���&�"��n���� b��!�F����B���ɈٴU�3抁��W��@�������W��]�f #�q��B����1�	e��{3ϟƒ�o���x��Q�)�ʍ�Ȏq��}`����}\��7�;N���g�n�����M�H����z67��)�| ���-L�*�^f,^�/���ε�h����!� yy��s
o� � �.�����z�g�����y���r9xET"Gi������)P�W�����2@Ы���\��Wծ��M�`�4��o�c��sߎ��t���_�Y���W׍Ӯ�eL�R
~���0���i"�l�������@�?	&�V0���l��tahx#��m�"DS_�T�S��Yݪ��xZ�u���~!��$##j�@a�G���R�%L�o���\ڇ)�FbK�ÎFc��qM�� �s���>@	,��Ăh�=ԙ3�}H�J\[���k������*^�֋���d�q]\��vW@�m%��k�6�7����7��e�cy
��Np��ŉ����9��R��j�����(��-������dA�]���|�KX��
�U���J��[򁶝v�����$�Iv}©�

���,:ޛ�t��SErCw��a����ӂ�u�N��f�=�Rؽ�cZYR�^�� h�����ٛ@N"�c�-	�0���/Y�磭<����i�I"�h1j�Ÿ��=�j�|�����_|k?$��F=КO�r����0k�7_�sD�]�f(�glx	q*�d��qF&Iؠ�����Pոc�Tڐ��t8֝��#��W��u+�)�QN�`4E�1W'��wf�=Cs�S�1#;B����7��H� zX��ml �Ҋc��7�nK�@+���:�%�}�#���K(K��!J���UR���c�m���xe�g�O���!)U�	M�ʆ�8R�J�鹿��e߶��>�g�V�����څ!��b�$γ�l8�2�:�ҵ�үztݴ��}��J����_�VQǐ�SS��c�_��-~�krd��vf�`��B�
߮�pD<�@�_�f=�_PK�����޷�sH?�.�ђO�=�3CG�(�b[]�e .O_����n�D}c�|�˨H.�)&�fzMa$\{�DE��Ρ~�FZ)�Ay}kguU?�j�*3a�I9{�z�#2��/2'����l�_���{-��B�v)x�#������~�bk�2?�j4-������qE7OJOE��J_v��=	Ց@��.pC8���G]�cX*���ױ��RE�6��V�тMM�1�%�A%Of���Jd����=�[!j�CA��7�1��畬�^|�T�z�LT��m0�Au���+ab��_�:�8�e1�fp,OA�a�NO�����4�zg��k)��{��7���G�E���-\�=�Ҋ��ͩ�������&�P.O|�F�_7��Dm
u�6ּ���W�]6�8�k �I���u�n9��]_R3�L1?\��m�j��~��t�?�xu�����`S{�N{'xNh�)��:��x���e��]i2R,4�}^���.)Y|�!I�����҂�s�B|n���g�D[I�"�qO��{K�	��ho��~�ƕ�bM+V��p���AC����/�um���d	�c�;�ʺu�=!9~:ܒ �������o��Xnbó#4Y�ʂC����[�F7�h0q���7/P/jEϷ4��LW�Q`��y�[K`V|_�ת��@��V�8�`��y��=Q�+�[�r������������=Mc�r��5й��2H���l�9�^�	oNuF�}~	x��ZT Yk�:�8�QW�	�w[k-O��y��WV3Wv\��B�Ԗ��$�1vFZ�W��:���葳�4,&�o�qGj��D���>Yk��Qr���b�mL�+��:�$�OJ7�Nӆӛ��ss����,��-��g�����T���u
�"��G����?e��m�?-FG��TJ���9E҈o.��Y�
bn�Q
 ��0�0n�C�?M��&
Kᡈ�� ��"��Q���N�
�(D:�8D8�':Kͻ"�H��� ��o]c�������xܲ�*dքx9V~Z���2t�k	I�͕?�u����>�(Ӭ8�c�sO4u�w9���ɢ@�p���ϯ'��*��8�� 9��� ���	���lM0a��2o����	����ED���Zj���:�@�aI��hB}���7n���1�5hF��Q�>�A>4 5���3:3z��ʦ�ÿ,ل*n�(gC�@�����zݞg�6���\��]z��G%��c3"���~F�`R8���s����j=M�8/�.N�]� �	<	�Z�W1���}�\���#��e� �`+�j�^�J�b#�.-T<>��zI弇w����ʻ��C˃����K���9y{Y�����������4���ڇ��)�\-��o�;gD7�*�FEo�Bϵ�'(��=e�`6y��	_Z��>pw"��7v։!�h6�w�����=|�t�7]џ�ZgyN[�l�^-��yܵ�T	�CQ�Xi���eh�
$�H�rdTVĶV	�k�`�:�;So'��Z�G�Xd�����c`�M/9颌�����q,~���bJ���%q-��|u~�y�8|#�UV���͕.IT1�Gb�:�Ya���f��ׂk�[��lv[~V<	��#�(`�.L[�f
8+Nt�BA6��|~��p�RO��ɹ�� ���mH��g���r�zӅ���`>��n��X.�`���f���L��HX{g%�H[+�>'�ۛ9˧����&䓼�������^b�(K�iZ�c�ȽS�hG�)�XU^R�ݭT���	�7���
��6
?�3���[�@��?64���?��5Inȇτ%�R��0D�c�%צhP�1V���3Ē�/W'�x4e�G�U�mB�8[�%qd�^8/鮐��9E_q��4��o�>#��z�b�'�;�J��� ��p�x^�>p����j�Aj�C�X��4��k����̵N
��y��l;��I_aV͹�"��f�(��EӢJ���6��cLuE|Q,�4T�u��Z1[���I&XVX��D�w�Y�OqV�V�̱7��XWs�"�l!�[��V�s�3�M��7���ȩ��.���
L}6s�r��`�}ս�v"�T�����H;�=�T'�F���|Gr����D��Ӄ������\P=�k��b󓯌�G"�K!~]�1oɔjU�1�HI��>�K���kLh��!�����Y!Rq4� ��|֊��U�!�$�֪>1Ґl���F����ax�!R���WO�P����S��hq��뽨��d8�9��m���Rb���i�&�:.�o:P���2��o�Ϛ_�)�7U�=�SƄ9�pye�S�����^Y)"�O��
�̡n��><��P������_��=�9�aUImu*ާ3��:ǵC3_�]�ܧ`�:��BT������Ax'Rh�>+���<_��X�t��}Ch��o!bo h/�(}ם�5�L%cC˒�l%�2U?aWv:���@}#:=r�o�'M^��g��0�Xa��6�*6%T�ߠ��f�Q�vj~�pڀ����Xpr�^�ö[�!;>�=<p��,D^�]iߨ���iT����&�s�T�ޡރ�`�&L��!�-#1ճl�o�G��so�5�U�l��L_�ފa���|?���ɠ��X�M�V �B4���懘�g�gb�x�&�e�I֫j�x�t:$V�9^�.b� uocJ�ܿ�Ʀ�!a|�#�ڐ��o���f�<��ݑZ��L�X�=����S����e�ɧP
nQ/skT�R��;2�LG��n��*�wwvI�
e�h~?7c\0�������k
�͵�7�S��$��zı���n�"��p�H���7�̩j����Ҟ�����y��~E�m���ph9K�r��7�~�V�/o	�
�����=A��)?�W�F�x�J��NX4��Y���<���Ѯg�G({��k���W,RR�#��Y����7���(A���-��WX�V���{v�0�;g��!������f�fB�?`V)D��j,���*���ވSar�'��8�A2����!�-�Cio�+>~k[n֯�3�6^%�吓�ńO��y�0���󮄐�#%�(���Wq�s&p#9�j<�"������R\%7��G�H�0�H��]�J
+��B��y�d������p��b�L��mDL��,<�Ʌ挛��y��*x�ܹr����gм�x��+�>w�Hˎ��8mM>k`1����K/���1�Us��tu�,��g��JZ�t>y;}l��dJ���o[��i�������p�)H��������D�H���i�G��{ ��+��A�\��>�,j�Wr�۵B�� Ѹ�9>�z�:�\��f�Q��p�
Y��Ń���a�s�c��s�[�d�+٭"aF����K!�t��M���ﹷ��\W��,lf^�-������8ܩ�Z�ӕ&3W15���h�3*��)9�ɦәX(��f�s1��1�`E��r?9�/��fb7��0W�6{�1�D�uP5��e�G�I�H�M�N�T�����]Ƹ���=m{'�h��)fQȥ����t�]�*!<mn�U�0�L������u�N���i3C��X���Mue.�˴G߹��C_Əxѥ��.VE��-g��hΝk�H�ˍ�����&����!>S���.���|�q|��|4 m��a���eÖ���xix��J�:ڠ(]�w��G4��׃��@�S�9}!������RM�G��͎*t1[�|Ү��f-�ߟ�@��I�v�02-�g3Se�
�{�n��d��X{��Ǹ�Ð[�L���V���T�{�=O�'N��?�l��Q�lS`�}#ؕ��?Mǧ�#�X{�C�ߋ� ]��pF��|��)��+��9a["���+��B�`�q4L\/*��z'��aëO�l�����;���gW �_��=��-w֘�<Tw�o�F�g˼{����<�$�&��4��ڜið�	�V�)b���l�L�c=tf�D�d�AZ��sꡗ�R����2�i�g��+��3��;�N��+�ȑҝ��{�����"��ކ��X6a�6
�������`Ϳ �q�4E�'Q�DL����L��o�w��wսu���۩�B��M�N���q�q��<�����h�T��V���
�%Cg(-�;�<:6�}�˖(�@��Z���f:�$J���R)D�#�1���s����T��*��jd����x���f�Pqa����gg_�?���p�g7��_��A6�F���,l�e�t����uk�5���T-͢ �Ď8�Fۯ�2$x������ʵ��f�]��Km>v#��↫�բ:�#*�N=�A�m򐙻m\�C�l����Mcl!&�iMEa�s��s5oa)d������x�֓Z=2�فl[�W\��3/� ;�/XԞ�8�tT�W�7P�5@Ќb�����>�e�B�߉�Y�tĄ��펷6���6ҟ�.s+��}+����d���@��jo=��`��������(���c��z��1�Qx�u�O"�����O� ���bP��e����͸��Uh��)xe'Rz��1���DuO/��D�[S!�i;Bx���Nj�[��T�;t/�{��/J8i��@��&��lHd_xB� )�){�m�E����I��a�t��#H�1~F����{s�	?����&�55r�������X"�#���� ��>�	� 1 w���	t���]�3�	Y:EP�>~��u��z�L�A.�+�Уhg�kړgՔޕM�b���@����k�=��"���nv�?Rf�Ty��m-��T�@$��f�Z�w0v7���3�%�Q��(�)��t��}%��S����CګZ���!Vd0������za��xf�f2��+/�ގ�Z�
'J��z �9�&����𰏺�L9�4���?��īZdZV�ھ�%zUr:�9���߶I�7Ae��>_��l}����w>��K����
y�'FjPl<mIF�u�y��D��H�=n"c铒m������d�g��*����᳙�+��>XoD���7&�������(�R0&�L�g�K�*c���U�#dM��F��ۻ�|��-_��xJ���
���-�3N[Gf�iy^a�e!��#���ؔ_5M���풊������s�#e|�ک
�T�I��CK�� �8\hu��/ ��?��w,GTo�{ �[T��&���ݫ����\�KQ'�X��5�ff�q+��fЃ�=+��@��p����u�V.�����`�Cf\+&��|�L��2H��G.+���9ɍ;�v3����C�4���6&픋��{>`�AӉ "8���,�D�#�
��+׶�w�|���S� ��{I�zBoW�i􊭪��M�ݍD�Qtf�Ec��ρ��_��4�7ͤ|��~�;���pki!L�g����O�j��`��;a^dۢc�A6�^�a������OM(���Y�8J������uΊ��g�¼�G�́�V��|�K�o�=%� �u�>�8�>ˤ�sȱq�A�z4�v��=#\���|@(|$�����W�w���M��g18ڽa�Em�9:eQ�H$~�-�����G���^���G�=�H���ݦ���,}�!PzOF��A��ՙO�Z��D�L�x��{�B.�xƳv
(���]q�_@�ÓB�����B]�ZrD����EлP� Y���r� �:�Zs?|����怀�8�9���ڎ['5��J��[o��$�Jg��P��H"�K�nQ�ls^���Yʍc-�x���u�D3U�p���EpG��n��~8�o9�A��O˷4"�Z<1�����,��H��S�C҈+$��`�@�g0��-B���D¨�Z�r����ȾT@v�+sTG�Z2l��' ,{�d��2;mRi�;ȼ�s��~g�C-�p�W|�䒇��D�c1����9{ԇ�X�U?�u5IZ#v%ޖ釶�
��7�{*������6�j��ζ`���EH{�Kf���Á��� a����U��%���Q�^��~��AM� ׌�T�;M-l���;�}{��/���M 6��+Cgm��c���YN��B��2��?J�Ͷϗ��P���甕�6����N�l��c�W!�O~�6�d߁���9|!N���S��kI/D�9�p��A�̅�@E(���y�4y���t�<�I$�_u�o�O^t������4P���*��~�:��k�/�/O�#~<H��v�3F)���1��H"<p�]3���	�i�[@��5�Z9��bDJٞ?`��Q�H�Z����H����YE_���'�8��p)��U]_��9�5��_l�'7}0�R�('�{3�H���Nz�P-�i�k�������c\��rc[��*H�$�M�eLZp�N��m��Dc�d�Ga�̹�9�{WY�`�E�w�hd���5*�3�J��O1{�#a x��"fZ%�#���-pCڱ�?���c�x��W����.�XU�4�������x�	� x����	w�J�,��x�H	����i
)
Y�n9�����Q�Vm?Yˇl�̴������N�aT�/*gyʚ��Q�hL*�{�$���׷�3	�p�ĢS]tU'��}_Q�/6��Z�����q��U#�ɗ����9�m,k�:yk�	�U߼ CY�I>1n��!4��Z�&0[�:2�Q��*E 'T\M�23&*4����IzUp�"�@�g�<�1�ذ���dtsmԭ� Bt�v�	����H��Z�)��)��栶Y\��~�l���`����&F�;*���o��x�(���A�����Iy�v&>Uʧ��u��,��RR�����������f^,hV"^]6�Th�p�7"ȝ���'���l�%$�
Ԟ\�6�<ƚ�݌�t���,}�>X/��Mfco��7�����a��Ԛﲵ��z{�ю=��;��Z�dqI�6�x�F>_���V;>��T�w�Lٖ�di�ę"��`eh���[p㭤�e�=�OP���r���<Z$;`ܮ�G����9m��V?ڄ�0Go#��v�UKK���9�5����5^>�<pMkV�mw�n�h8<	0�A�=1�7V]�(���w�3$w9�gG����L�L��jV�;h_��V�77յ�|!���M{����:,cI.%�R�X�65o 8LH$���xМ�M��u=�w���E5����J'�-�#�F���=<D�R�-ia; �L���)QK���(�������4����8��tR��6@D4 �%Ͷhf�y�߁������q�+d���	D�ϦͯNB��[Huz�.O��vؼ���H�75�?���w����L5Q�π��d����D��2����u,����\pH�!�^0�J\����d^z	����7�ڌ<;�ܥv����z�"�3�EaȠx�@8J��:��c�)�C�?�i�����E���ah��b.���;O�W��+�0�q~��C��5aT'��e���ԟ!bE�� s!طO��֬o��CB$����୔�P�$�H�s!�m�H浒t1�D���(��?�C��DP^Y�+�m>��xE���*'V��Z3��1��h�&4�y��>�9��Q�7,�>��a����F�JT���P��J��՘��k���Dʗ�
��c2S0�Я�B�̷kU3���|P�Qund�mv6v��y+��I�2�ɟb^f�BE��|�!x�3��6h�P.[I� Qb&��W��^������F�)��}�;	h�\j���n�9������ńK��n*�[^[ܪ�)���uj��t鮢��^��=��m��ЪA���×��>1�abC�Q�Tx�?�ZU�1�"mg�ɍ�1rTsu�UN���� 5�;�����>��R.��o�i�{]�1G�y�b5��`*ALO���O��3u�ް��}��U^E|��g�2jm��D�"O{��WR�
<My�  (~w؟$r��B��ʽG��V����	j��_Ծ��J�)�,+A��J�f)��?c��=�4��Y/��*��'����3�v���h木��d�҉��
�Ef<��\��cB���#a��C?�^�2U}����*, h?�x�����+��E�Dz�H�Ѱ?k �d�� ���Z����,��"�Z��������_���"E�r�~�Ƌ�`EAW{i�H�rV�a�Av���pM�8�(�b֔���}B�pL���R�4?�g2$��`�Н�[(��g!��w���n�y�737�=�"tOW1���,d|��diTx��$g�˫6��N��宓��CO3=T�[B+�M"䘯����l�5�)�OWǦe�%	���������/����<��. t<�.x���0�%��� �/1�P����"�����'L�Hs&�C�fmK�a�l��A����v����1"_nS�%6���~2]��
b���*�����>�-zS�ifi���~��4�B�[�a�% ��E^����I�$���/7�A��@���1ruw��������"@�����S�'���f���M�h���hϜ-B���«&�{ѧ!�����v+G��Y���6�b}ϙq^�B��fu�mHq��w=[�Ӎ��wA� ��}�D�T�!�Џ||A6OЖ�f��� Ǎ�T�CJ��j������Y��,X��X*���p8�Qz=`��id����X���ą�&W:��s�`���3z��m��R��ʲ�߾��`�5���w4fyX:KL�zm���_s���� ���[��x�%j�(~B-x֦zm���&��u�FB���,F�Ӂ��R����ݤ����Hl&�֓�ct���qS"}�][��Tsŷo)G|J@$����A�n��p�t/�����ܔO�e�z4��Y1�����姊�u�6Җ�cn�| hd�ů
��Än?�8+ �:�s	�e�T���"hLǭd4��~8.-ҩ5I�4q�쨙k�k�2H���b��GU�~3�����hi�ݐ�ụ)y�P���(���Ɨ�}�kP�=旸c�؎N��U7g|/��gl�'��k�J9��2�K���Z�@}hTI�XC$�,�X6(��\���JwuGPjh�y���	*�v^ϟ4�Ĩ=mI�1�C�E^�0�UHS�_i�f1�ĚW�C���9Ս�ʣ��6����������ZυǑt�3��uP6P9�L�	n�}���=�������@�چh��$<�R^7��������ӑ�8�Eo��\��-�$4
c�].���@�JL����+"�) ��7��F����mO7���C���L���	�b*Eyd�m`�{ot"g�ٰ�Ui!ύ��5�l���Q>R4d�0�}�:=��N?��c=�xz����cӭ��p��Aǌ��(��sh�8̘���Q,�4w%v��v��u�W>t��Qۚ�y���(�@��wjL�#Bt�#��p$���VS*�Mï�7�����x�1A�q�OjEXQ���*�XM�aAo��pa�:®^��7��R��5�K�"�0���~��Nw�u��x�~xj|�˙�X�%��%# �Q]}R$�4�w�.Â�͑�_��Z�h�����ؔ�����hf|���@�;�KTg��]_���^�؛ĜK� eK�b$��$\�û���\K�����[��<�6�j%tSc���\�ʿ��Q��s1�2�é
C�(������������EH6�T��[��O�$�iz�2��ߥg��5B<c��l�K���G�E)WH�?Ж�'fPC�������W��Y������	a1�~��+P��@���[k=�q��W�k�cE�;�^���1j��E�*�����Y�蓕�f���]�M}���<+������>Bv�|�Q9��=�~5�1�����ng!5��͌��pE�Ķo.�<����:���*�7W���"�x���#*9���Q��l �c7ݙފ$ѩD����Y�"��,�}��N�\D�7�����/ȟ�߂@,��/�L?�
��3k������1�Ꮧߺ��8�}���/-n@�r�A��5V�/�]��&�9�$p�"�ZC�D�~��Pi�M,˞D��"s�$n�p�5�MY>��x�%w��|�J����$�뼦k�˂)���_��W�CדA֝������Րh�a>�ӻֈ*tA�YLÎ�a�ĦΎ��m�R&��m�]���ڶ`ԝR������Ɛ��5f��^�0C���zy󛍠MF�S��0�Dh~�!x5��b^j��Sb�;�� i1��d|�Y8��96Sז~&���J��W#qg8��B��߇��Ċ��3�o���x���t��.���%E�eJ�ú����m���x��%�g�9�F��{�~���5��j���5�O�.PU�����A�T��j��CF������,b��?��)����H�H��S�)R�t�Db�1�&NƲ�%�J������1��}+��iA���:5S���1��7Am�+%5��A��JI�>98����_�;�r���Zən7��z��4���lN��GJ�����^��ݺ2�,����-�q����������/H�s���s.�}����oN�Ce~X&�GQ�����Ú2�(�7�t��-$�*�������Ma��%ے�����sU��E��6,�߰��\�x}Y�*�$�v����L��UıWwfX㠭��wH-�AIh#Љ����(�0�o1�%+�b���+S�S=�E�9Y��r��e�CE�}GI!��|�-���w�y1r����N>|)����U*�͙D[8T�a�}�qr�6j����(>*�{���_w{ҥ_�b}�3)����i�f#^Ԑ�C%�V��]r*RE�!pw�̡diT�ee�Rv�]��a~��X6�X���E����}nZ�nƟ��dPx��d��e���@�q����ݚg�JhV|	?��(�E�m���V�Y=<�(^<$w�ʌ�h���b�`��H교��y���V�^�h_���.t1�Ie�k�Z���H��E�ˠ��A'/�˞iɨJ�?cp뻊����轵lڡ�Uc�ʛ$7 �S�#��K#�Vm%ߣ�w��-t�δ��[*^�����ė���W�A�&� ���x�?����J	K�Lcֻ�n�r�I]���AR�L�\�(�^~Su�l��<<"��)k��k�p����c�A�cCU`3�x_-���WЋ*b:��lnp�a+h�Sa8`%���Y��Xb���%^��MK�Uh�Gn�F�l�Led�������! !w/��F�sX@y��˞:�;��jۑ僵Uw� �j.r%�F��T�w������ȗ��G������ ]$	1�:dkorey��z_�RI����H�)�'��uD�@�u���ͱ5��%@/t���n�x/�ի.F5�썯��pTu��G����D?�7��Ի4�.~Ĳ��h�W������	�g~\ce� ��3S��<��<��0dD^��fq���
��n7�)�I��+�5ݱ��NOi�wR��zʛ@��ٗ�&�eK��م�P�<�]֬�����yǭ�>���F� .^��$�h�;~�j0��\��'�Ѱf6��Q����l�F��R\�qd�.����g��u-m}n��fÄ6$f ��CW}X��UB�;O����3�����I(0'G;�[���\�5KC�^z����*�b&�s��/7����+�����^l�G=��R�f���(T6�@�'L)V��W<���Tܝ/o%��R�b8�zi���$"K�����g7\��������?#z�����׳��c�R����z/�&����|�$���C݈e?�,�
�4!�G;�B�>@d��<n�d٠*�*Љ�O���`�����J(�> G�]��4Ǘm0���^΢�u�}S4�筁�WhHW��Ń��I[�G�h�.
	�Ϙ�6�1��
ܪ�L�C�8$<�'n�!�@�ѱ��⇇ݦN�����8����4�Vtb��(�W�Yr�*��:�"qm�@�/�"]�<%�9�'�Saq��3ze4c ��H�&�F���-���y��2Ln��� F�>�m�[�ۚ؇~}2��~x���t������"�^�_#vrǝgشt���̲#��$hq��ggxw���}�t�4��Ck!�DfK0@��K}�a-QVD(j� �:�kҕ؅�PY�"3�=x�c"�|�a`H8(KZ]�����iǋ�,��F�V�@O�nS�{?-�1.?����2Q�'��罚�)ts
���bG�Y��N@� R~/�6M�n��!�;[,|24�����V�9���x��E��9���<�$'��d�����\ܮ�ܴ��rB�}Y����G0�P�&� ��f+��vFg��Ɋ�>���˃>#��˾�:�T�����x@=d��Ke�2�Ƃ,��S�W�]d���I�٫9E�	�览Su�2��*H���w���؟9R�����\j�MBh�m;K���@7�<�,a��JسCr�3\̛^~յd����$�M�6X��1?����-���������e:	��z����+*)�����)�|c6� ��.��J��m����5����[\UV���x���be��f&����(@X���\�� �&!�j�M����U��3����^h;�x�ا��:NWH{��|[����W�Q����P���<fYb��nu�"�
��F �Ɖϊ��[�M<G�'fqW�(�#��#M�!���%�_Y+.�?60�23��Ǡ(T�?ݪ����=��װ��(dLI��e�XA*WI�9�Q�2:�n���b8�+]��c1��blS��][�D�O$���)�˼ٕ��7P܇)�8���?��Gg`#�p�#�ks��� ��}�)}y����ň�t�����9=����km��@�Đ��x��%<�|S�~kv��{�5��&M�L����B�f�AP1�)�G!��Lo�5�V��9g|�Yy+W��]t^��$5�闿�BR�-B"j ���ґ{u��m
�������1�:xi ��(|�;٤��G�{��?Bh���w,��g�o{-�1��Ye�I�����Z� Ͷ?�����y�&� ͙K9v�I���3�>���Ԁ� ��[Z�mE��D8�����>��?�Mx-�3�%��B�$�hs%�Hl@�����5Y��qm ?�z���I�P���4	���X/������ʜ�$;��o?&�h�^M�΄��G��S%"o�|��ͨ��^@AP�ߥ tO��IE����E�,C�u��Yց�\=�b~l=��vGu� �'/y�,�b��7�x?��j��͹P�3z�������Yο�QZ�󘵜'��:����K�X��mM�W݃��Ǖ��N�ϋ���4&�ә#u8O q�I����8��CV,M>������T>.�F$U�2���w�>���VP��t��>�s��s��P/I�C�0N[~	�^DٹaV�^;���8��-�[�|b��ߠ3���?7��-E�1�ŝ�x�햝Sr��a��&�!?n����)�y��,zR�e�� ���k`q�����I3[-��<�,�t�7��םe�H��+��ͅ���/(w�dSp�V�NT��nI�j�k�
�9��v^x�d:˵R�n�D��Lb�������ZA�P��i�}��"l�?8�W��a06as�D'���J�,;���(��H��Fip���K�f�3���"��!������$Ąx0�����3�L:�)#�Mb���"7�W�na��)�����z��B�!�iј ��{�T��\����'wl�]A/-�f���.�U��pd����� ��AØ}�O�w6w^@ꌅ���q�Ox����].~*��} �a�~P�q,�Kw7�������INB"PZ������x���t�t<
��[���K��k�p��b-Ќ��>�	�h[rG��F�Z�����I�����I��%�q��v�{��w��j��޾l���?l* 2�'������w���O6��Ox�:>|����  _����ԧ�{��$��7�ۍ�����)4r��~nJ�m�Pvt��H����3�܃�򑴪h.���mЩ95�~�n`�����I#p��<�1aFȦ����a�7q�ncc�É���s�E��o�iO��؝�7���b��GR��st�������1��B]�НI����p�|�R�'x�T|�!a�v^�U{g��WN#3p�C?�����pu6��s.�"�B�qVŰz�0��zZ�h+�'C�B��2=��z;�����k����S����"dz���ԗ�,0|��� )��yM�%��U�Whc;ՉtM&v`P���Uu�y�ﹲ?l=ۮ��~���P�)�	��g�<tE�b�B7�n���������a�ə,���8�ao��'�s�{�v+K�"�ጜ �E��'�_ ��1�zS��E+V�g����O�'�PJ2�X����R3������C	�a��"ady�'c
���|3Dc'��2�t5Aӏ����5��\<H>�b�(v3r�	������s��f��N�.�q1�p���4� ����B�E^~�j���j�����O-��D@q8a��!�;#Y��Q��P��#��)U����F����������.�x��$��;8�Ĭ��S\N����C��N���\�y-�K��)�T�i��N7�܂Z�n���t-�5��AO�zG���.���5�7�&#���b$'<�Ǿ�c9=|�ށ���9�ΘbH�d^�34!&k�o�k"3v����"�N#�Ւ=�×��D���D�6$��/��G�*��Z������mՑ 	'4NF^��8���G��Y)k����wt,= |��"�-���X�k�[�*V:y<h&���A'��7�Y�;���\$&��|��p]*	sN̊Ry���nM�{��i+�պ�KطC�nx�Ng��|A-hs4?�0?���������<휸[���s������Mj�_�43�glO���c��W7�(7|%:G7\}�]P�۽P�~V���V>]2��l\��, ��ϳF×tt�>�I}�7���q�if�9�Mfh�sg�`2ߊg|g�&���9D������*�Z�9�I��}N鱍	�[Lm�Fo��P&��S�&�Eh��9��hī84��1*����_lԾ��X���
��+�*�*���J�XlU����W׊��j�t���ȼ�u��,j�cp����	#�m91�k��13g���Ó��3��>�I���hѭ�I>�#U�6��0M�:� �4���o�
]UВ�Ne�-�~L��M;�;�{@�M���(D���� eOW�����e7�gp���.��L���*u��L�����7���̴K�c 7'v���3��&�{A�E�P=�����Ona���%Ӽ�s���z1��w���7jE7Z"�'��$��f������3��R���&0<Fe* �ŗ�l�JIn�7GH��d;s<;��.dFX��쨶:�o�f������ƥ~��m2�~������e�A�Y��'l��96L�$��D���S=�A�&�^�-�R����ӝ#�T)4]c2��O�`	����o����o��;c�)�;��8�uפU�K���E��%�O��8Z�̛.:��FO|���̦�S����-K�=.l��x�n��fB�$*���+=UU�C�C���EP��IL\�`�����Y<��������fRݼ�46�O���s@e_U-��"�!u�~"����'!!>"�ID;�J���^�#�ڛ�W�L�˩*�b�*�'3R����ū��A��J�����شH{Ll�
�ߑ�K��0Xv�mی����ʡ+��{WJZWXd�� �x\�Hd�����j'�u]Y�,>��@�m��o �:� )��:f:p�Ԝ(w�l���O�>"H��.SY^6�(<�Q�J^�O/q&t�	��*��{�� 3�U��x7���D���΢	H�����p� =b�t�!ʮI�Nhn�pl�����_�<Id�؝�?��n]#����Q7eH>[��v�'-���t�BVŖ�4:D���9�]B:*q=
�衛N?]��#Y+*��.�}�%N������kA��w��%Ҭ�7ޚ�_En?���KAKuܲ��<�@0YK��C@�Y�M�����n�s!��v^=�_x��S��F�m�����Tn!%>g	�\��Z���2��w>�ܲN�g����N�J��ޢ�s�%��B���
���\;�'��d?��zW����:�Z�)⯖�[�Q���w�l��^'q+�h�.:"�T���̕<�W+~����4��D[��+��G�0�[��\(p��F���`[�ɹ��WN������lT!�V��+��q��.-C�16�{ �萷��y�x��-��x~�_q�b��ҽk/Y�uH�����HkYvC#LR���X�����iR�F���+�;��h�'���n�1�{FX��D���=��ā��z���͟]#�ݑ0���C�����[Z[,����O,<j�{���:7�V�����a+,=�8z�KC�a��R����7h�"K�&�t^v6��kY5U:������j66�T*�Mz�i�qL]8�mQ�Xf68
>�|c�n z�;o�������ŷN�`�;UoT_�h%7a�:����h�U�!��hFj�+K��V�1^;�a�Io��$N�e#J&���64t�2�uX���=s�@��PKO�`|-&
�~��j�8SHg��z��甚��9��HJ_ mϿ�H�|�s�w�VL����S�va�2�fCN�e���Y���G\�2���490���Cg��x�o�I��B���0�)���>�P;��D��a�D�xؾ�`����g��=�l���)[d�@^����z�E�����-6��ꂑ�I�9�	��ٱ�k�����&��E'(#N5��D�0.�G��2�AͰ}ցPl� "���c�T�"��U�K�~wtf����H!̷g���u��/��5�R=|�~�An ���;6��&����@��1�ᄛY�Yq��\CĈ�SY�v^�ڗF����F��y��"E�X@����^[F�P���LX�W}�X+1���;�������"Ʒfx�����@�!�L�fq�<��-!��s�[�"���;;�f��^T�UHE��Aԉ���;�%-�	``,6�EK�}��)n����U��곯a�_�l�\�*��Yw���)y��z�d�����&((�w�#�տ)/�k��(yt��n�I�v����~�IC���ͦF��U�N��n���I�U�d���J�M�Cc����(�]�v_��np��ʦk�M ���RI.�A�C��N�M�5���́��n�~w���'��8C�١^����j���Qk���i�0��m�!B�+1�H��N?*�����<$f� ���2Sq�wr=��%���.�?�g�|�/�FM?�b%����Y�#�ώU?�5p�ƹӶ��G��Υ{>�VDy�.�M-w��
���wEӯ�T٭̽�ǭ7���5:�!����(��w)W��Ծ�1Tos@wď���*V:�%?��U�z�"���E Jѓ����+h9&$�%Մ�@Y��Z�Ѷc�ᓑ����~�#���?&�����(�͝<�z߁��8�]Cv�|(��y�^�Iq;������[1�r\͠��s�H�З��"[��a�3�\Wh�~DIC՚#Q�m'��R�b=:�LP�O��0P$?3v�4=<���L�$��k��.����6����<O��/�f���Mg�En3S %l�:����q��4ç�b�.�o}�^���"'4���4ܩ�M5@8���,(;JpF�Si_$�e?���6�ɳ�H.{��a�Y�q�C�-/�sp2(��|�d��0�Ό����a���/A��)�l�g}$��=h Ɣ�<rbsg�9oZC��m�M�`�ҭs����eY�������J���uTc�f%v�i�Ҝ��;f���١M��i!?��)am��D�6lp�����yđ9-�и�d��u�X�̭(��)���WM`/��OA-�D�̘�]�2ϩM�)�����h|�~�[9٭?� I�P9epf�SD�2���+�����o.Fs��v����hd"��7��p'H(O��L�X��z����� Ńha�H���9��p�8Z��j{	�'��7G!r*�0As"�z�oh�<Io�C`�P�ɓp_V*��)�6������^!֒*��o5�RN��}�Ë{����N��gX�ʺk �-�u(�"�t�:�!�<"������|��4[CkP�r2�ɰ\˃��뎲 ߸�>�`���O�����!@_�[��{_蠞ۼ~��Ƕt��.����?И�M0��aTH�{<���VD*%g16�e��x��'��BH_����?ة�$���#t�G��o��ZA���Bu�d�6�Q
�����;wI,A��w�!��i_zKV]��o���9�9&���z�LlL޴�TM��
t��_��})����t���4��{�j����_b�*��x��81\�1�P�H�Ϩ��Đ��*�*z����
�v�{?��y�aD��*z�� 
�/���TS�"���|�IqnN յBkV��T�y�K��؁V�90��_A� �MDu��J����,���S��aKB����?p7�GNP,��v<�`��%�3~�����וVi$)�ӯCQ����u�]�ru��(h��$p�9:�V$���/�S��>p�!���̪��_٥�z-#��5�ǡ��R�K�S<T�yK1{�˰���p����L��H�l���dtە�)4Y&X��U��d������wŠ���K@����eNh����X5<�
�P�I��h!��1`Y��b�ŀS+�IZ<����Hº��Q�}�ףV�t#<�[�{���ݳ�/��N��À\x.�Od%�p��.��B�ٯ������@���!re1ypsA����w��Г=�o�?�0�Z�tՊ_K�,����#L���%bP�q���iϥОs�w���:8�������~�>q5��3�m�{BpvRE�A�9�JM߭��T;�QJY`r�lr�����lY ����Ы�l�����Dɗ�<��8�]��~o��Ȅ'	�B�%���Z`��bT����Z$ ��c��7��.}Aʭ�2��,=��i��E	u	IA��iv�	{%����4����h���;J!�ȫ�Ut� Ü�հ��0Z�B������VP3d/͚dt}�4x��^5[�d�|�5O)�o3�!&c�腺1ގV�H�o��M���o���6L�N%�`��p����cў��Ǒ��yE$���$����b�q�Y���t�&p`�3�Ϥﴤ�0��3���z�<3�v���	����N-/>Ck���e51M��
�HH���m�7���~�O�%++��F��A�<a�#�Z9aZ}j/Sm��:�
�<���l�e�}�m�Wٺjɚ�O���/����������"����:�6�k�U���������P�(ؒ*�6k�I�3m�e� �Մ;�/���b�����}���ad f���5.��)�H�3����~�UB?h�Ş'-�֪¤�nI���3���2U��t��T�N��6��bW�i�r� ����Q}�ɛx�:}_p��hh���qؿ+���I���M�DWf�➍�hK0�_�7���kW����+���I{K9�����%ƾjY�j�$���
�<v �	��It{oW�)���V��(	�_SeWlY�M�!��="����JJ%���.�:�xR�6h�E����ƹ��P��:���q��~v�'Z֌k����2Pjl�?b���_\����zr�6�?�jC�	bm��1�~v�6b������ͧL��&ה�@n\
�D�K���ii �
��I�����%=d�C�n��V;,���I�c,�OX�yQY	JO�VW�nͺƩA��[�l��!*c+|bt���%W"#]%��a[�#VZ�����`+�wpV��AF��P@`����/�ٿi|Fف�ʪ���B�OI�9IK�u��O�Hẻcvi�#�<��wn {0j*�|~�Y=j$	��η
�IQ�fQ|S���;���c]�1v�0����,P�Ol��v�]�D���m߁0ۺ�!�n�<�]�r>0GB @�u�pz��J�aV�L��ܟ�|�y��~
�#�:��Fʍ7h#�k�����vX)Ōy;��s`�,�ӿ؂?ZZf�r��yd/�A2ZtA�=+H�O��txq
���$t02Bd��;a�l�t�!KK��7�؂���֧��K�fwI�q��Fws��n������|%������I)Lp�F�@�|��k<+��N��|�������n_E����jX������e�R�(��*��-���$$��8����<�|�&jt.˯�FW�r�]�����y�/�s��X=�MQc1f7��M��	~L�R�5D
�b��;
u~��4��4�]9p
nF��g]��	ݐKΡ�$J^|e��V(젠���5��]c�~�1HE%��6����t�(�(�k���)�͸�+�wb�Z�V���s?1�^KD2�"��#��nV�ICG
%��Sm+^�l�H"Ծ��s��8{���Ve��d��K
z�ϴ�������m��Q)=!���\@�v���i�hř9�w/��U��$��-]�t[<��N�0��\zb�iS��ǤO��0�>L�|˻`�Vq�MD@KtЬ�y33��M��;VތO�?#����v���5}��*Ru�`�7�����v>�x��V6<� ���{yŝ_�.���~#X��ɹ⌤�Z��|g��4�z�	�ENݼ7	�m����X)��s�kv�Q���+�f�=�,��M��"6�@D�5�����p���%[��p����wV�7.��Ϭ`}�U�nvr��h�)��O�F���\EW��+�d:�;]�z>�D)�^T��Ŕ(�y0n�&j���l���:��X�U�X�JN#����ْ�3�xYp�h_+ ��&9E����1�@��.ͬ�ܠ�\�iz��kV\�:�	��#���^.C���݊�gȦ��\���D��O ً�j�2oI3sf���3Ge�+��_��tO}�����Z�^���t,�>F��1o>�)�����C����8�3�>Oځ9~��_���VvgS(�˱-2����O��`��xߧuo��iDv'��p���Jg��Qc��$��l�S�(	��bu��:��h��DR?���N�ݤ�S���X���Ӥ6+����1������ʇЁ�>n�9��z�,�T3n��$�9��o�<���l!�8J�#P���+���EN�}		�5���E���m��������Z�j�.#�2P��Ѻ�H�vB,��Z�{�U�@Z>���w��_�.��J$�*��X��Қ|�P�����!���'H4����Z�U�zt��;��OU�w0�Bתzt��3��'=�� �����1�Y@ߨv��M%�*nA����>�5�*s�K2<���<�4�|��n���6~�h�:���J�Q�V�B�x3�(����b�Pb��j�
hNw�����N9��R#&ca�r��v�Y���]������C*F͋��tG+}1^��,��'�M'"	�iY�JP{4��>�����W�Fw�=�{���q] ڨn�m$�u�!����&̏��W(�X�:?�]�����j�U�͚@��ŷ��^��/�S��_raƒ-���CvԢS2C����R�	�<�yCw8�a�1ǉ�O�ό�+��W�p_�qK��YIv�g��r��Bw8��3Ju��f�OdFJ�w	R��Y�S0��U�g|S���Ob����!�Q��c3����v.���"�Ba'�$����P�z'�H�"�����5_Dw
��ҵ�9	X+���Z�y~N��ų5�P������BӞ���� ؐ-�Z�3�j4銎����ЈWw��`�!�Vs��@��reQ%�j��y�	�^��&t�!RsE�Ӱ�A��~Y�5�U~}�{(�+���N~�hI����oJvHȦVҵ,�S�o͢�f�FQg%�Z�Pӿ����J��.��v
�X��A���ZBb�A����#4�w��.yJ��B��V�F�iy��s�bvEzQI_dި�Ñ�?U����/�b�څSA$��G�ó�"F�y�VN{�;���/n=��$��ʳ;��1�z��m�'/|"�"?�RZ�1T���X��=��r���j�[�ߋbW�Zɴ���NCb��q��'VJ����^!C�=�	C�&�A0߉BP�S����z�ܻ���Ifq�v�w�p�в=�/rX�'��%ӯ�m`^�rg��4_�R6�u��>/N2���i�L�Y�r*̏d�
$�>*9ѭ���d՗^����,EHc��WyMFz��L�|L-(��7m\�7(>�7z�C��Pu=��2IWy���  *Z�C+����oN��Ҕ޴�U���K\���L�A��V�>�v���$2��ז�K�}B�6����9�\���<�`<H��An����C`x2R�z�a�@~Q/�����#�=�$K��� �8$�C��q����%T��6�$�
��qm�hX���n�c 뀎�	`F�MT�"�Ժ�d���6n��3��W�f1�Ȓ>�d�Ȱ�Z�$��g�ќ~�?҅�����8�c�ʯ�0�3*5_�Ŀ�r��ʤ���Rm� ��6�M6<�`� ��[����O,ԟ_1*�D'}竪���#�KU5$"f����t�WE�3�?�\!���8���;�(�é�CL�����X�ҷ r2v��?L$d�Y�>��%9rqw`j'�����/?(7�9�w�̈́��ZH���3Yj��J�����u=:��p�����ž~¨��Ĵk��2����x,	^;1ɪM[��8b�I�.֊)\n�)-�nQe��,dcQ:��G�kв�f~�6:���k��!���S�&)w�A��B.�i���_C=м��~7ΣI����R,.��4�N����?� �X���B�� �>Έ��{�ei��4N��$\�yB)��b$N�7 z���zK^�"�����@)�1�u��K�r̈�M�-ze��I*��-'��kg)�����A�ؾZ_C�N������B�� Z�k~���✶����Y���-��f�(�'+k�2q�q���Z�'���[��p��c�V�2@��!/A��1A�/��:�9�������cW���%�Z��#QC Jנ4��a�Ws�J����qݼ+:�K�ZA�Ҋ�3t �J�iD�)�W4(����8�R?���\s�%�m�|�F�t��u��K���b�VaY�*x��h���oDw�K!�I�.�D�_���D��K��e:ׄ��/jώT�Y�#\幸H8"8("�%�W���R�V�0ߟ������w�+©����ʮ\ט]�����&�����B<,������L��X b�y����`�ex�F�A��q�iR�Q����;�Ō{{ï�T���9�%uKW�,t*�/��MP��[�g.�F{�#�Z��8��KZ��ޤB����Dv7P��	`���q��~���k��n�zh[����K}(%���Sr!1������~�����N���ܨp1�7�
O\I��� 0��;���!��M�
��Ձ����.?��Ě��E�l��yY���Uf�b�gU�����$1���#���V⤵扊�!���9�c�V= �1gh/<s�e@F=6���P�es��,J��6��`�S�z�F����D�j<�q)�y��@�y-Ƞ�u��
�]#������2k-9��z�/I5vM_�rc���ӸE늓+&㣫�<�[��Hd{�U�E|,�V�?~^�?���M�!�)lF��RѠ��yw;���]B�s�WQ�9���2ݍ�"n��n-y�8���wx=����f��,|�������ۭ�ƪ����@���}��|��S�!�e�|�>�;��|�)M�l嚩���՚�	n��J��ra(nӘxcz�8w?�������o�*��b�2���)cPe��抭�ȸvimT ?�����z!ŸL�^(��#�^�s�zVR~l��_�7pJ�g@�;�:뽳�t�5-�B.��p�3������U=���v�+�[��T�[
�a�d}�c-�pz�V�O��JnݴH��Ro�����-"�u�U��<L��*H@�ϵ�KQ��J�n9�2c<�vx�!��?�Ƚj��8��;hбkF뼟v94�c���`�-�$?��X�)ؾٻT�Güφ�,�m{J�L�`�rSc����%�������?Uns����|p0��i�ip�if�7~$]����E�������>��g�C5Nd덍�� W`V��?`�������㮪��B/E�v���~sl4g�-��i�"�Dw�Z �a�����Zґ�0�V?by�2��Y}b6�S4�����K����f�|YT��@chH�;g�e0����4�G�Ζ������.POIb��b���bb3�i��w���E`~���^�C��-�:V��zk@	��ۃ���U���Ǵ��@S+ڡo�ߑ�Tv�ŤYV{I�Qo$�٫e��[Q�8
���w�m�
�Ha������S���O~�����-*�w���iB�O*�w�0Dc�b`�=%1,S�7��
��`���1�>T���N{y{lO�ا�!�e:#t��*�kF2r!���B�!P��cUP��ӴcB����F�Bc���9���~ ��]�Jdk�<��W�.�Ȣ:��{���_x��	�E�;&.H�ggaY��Z�Kum�Ee��0v�gު��tw���檥�`���
t�a���2�&�STQM��ni�k�g�3@U���-��Q�5�jNz5XA��ߞvD�}�G}�P����Y\m`k�T���T*�L��<ޞU�6m�ռ6��-����G�'��` fs�1��>�芿���l��.�7��e�
��G�iV�^ `k����Ĺ�����#�r,~jʵiߝ�N 2G!7�����g]R�/�G@����6���!����¶5����Pzgwa�(&ɵc�Y�uW������o��P�}�0A�|"'q���'l��i�R��q[�Q��Qu	�W�Pt)�T��\�K��[pON
�*���#�1`E��L<d�����פx�׏�}���HLo���;��^af.���%���IW�@�'k9��w-|T�?�u񺁟s��C7p��f�Z3n<H`tT��(
y7�l�|/�2��^�>|�$��6��1Xm���p���������
�3�p-������]�;;F�VJC����;�=�q��E\Y*�!��I���2!O/I���LgR��g�B{�4H�)0q	h�cˇ��o�.�*�����d3�X.q���nt��r���}!�W��p�8}���b�\n�h##�;��)�g@��<5�qG�ա�v]���^q��e�!B�zZ=����Ы{�:	|���v��/�j�P�IfU�~�wvг��D`�Ĭ��w�	e�å,���`����h$MW�ȭ.��/tUbLۭ�o&A����b6�?7"0Ep��fy'wK#^����%O��:4)M���򴫩g����+�:B�4��x4��;���&�u�V �_5-�c�g?��T1�e�����e~3x��M�lNF���L�b�B
�9n#F$�P'g�8:�Z�/�m�q9n^~1�k��,��5�`HN|���J<=4_�;9=�e���P�i�Ydz:��nRS~�O����d�����op���x�T�2[S/�@���b����_Y��u �I]�ow�\�C{���#8eӤ�{�y&pw��U��Af����}��)ӛ���Lޱ���� M��3�[��:�ə6�C�T�*UIz�܏��R~��<����ֈ/9�j�p��%����^�$�g��Y���XS�%���t@�/$j�&�6�.k�pX�]���'����HN�g�mfz�?_�V\b����I�핎���uY�2��\:��[�Y�kV��]�Bݬ�;�x�tH�8La�td/g�Ⱥ�Ny�ãYM����Y,W���ͪ�}9�\\��a)E�1����%s8�z��~/�%�[���'a��\�u���tF��r��-K?\N$|�]���;:d�����lЗE� Q{�I.Z�u�d�m�Q��YJ�JFd�����Y�]9T$��E�97�l��_jp�Sm.,#�D�@c`-)�S��E6{��ƿ#��q�z�I��	�zbfm�Z��ЄRB�̅%@M���A&�p���
�N�#�n����P�y�X�����V�l|�OF��Ǩ8R<�$�G[�M�U��J�N"�	|��%y4G�'�o�kd���[���k��r��p_��m�:r�.��v�UQf@;@��GH��m�eh�ѻ�)�pgMR�I�
6�Ϲ�P:%��h����.��n�*��WbV�y]�#b��zD��=F�4oh6�m��hy�r������q/�S)
1���F�!KXzFHp��=xg����䟽�<jͬ�H�f�`r~��_��S���gL�:rV긣�v4����6:���[�Y*c�zٸN��	e�L�84!�xc.�c��������Bz�;h>?�v`��(oI%���,������ڼ���c���zb�p��=@D/��p9����`,�ZVN����v~f�;A;��l8f��T)�K�k%C�[�E&�����(1��#����������C�������k�<�R G*"��ʶ��#3���a�`�"X�,;�wY����U����ݶe�EU�I��o��k�C�ϫn�P�rF�Z0v<�s�Y��6�Kbp�X�R�#]°��Z��	8�dS�8�A��x4���[V1'�����6�Ѿ�*�D�~�uV��2���PQ�����H)�$�c�m�*$�#�1��+�M���wu��bg�o�%B�G[b��F�b�@�$om����'yqtc����t嚤7�� 0���+�0�G���q0ǳ���ZƠ���-ʥ�.دf�f��ok���	X'���+;�H)��J���D��
d�%���ḧ��g�,�x6u|l[OzΑV5�8��S�E����2����N�z?5h������T�����_�&��bo�W�7� f3@����~���.�3ᣝ����6l.�[��ݠyo�
 ׄyD�T�ܪyd�T`��M��!���/d�*���cafmmȉ����hR"*Sb���Be¡��#�a��NHo�O��U��eU��O��O����������i�x2���Ntq���y�2�N,�m�±eWd��\[c6�E��z���}�r%8��?F������v���g/���/P��[{�)�B�N�#|�{K�'0���˩���qc4�T�2�vXM�'ʢ�J�!&����I�4�����D��yy�Y���]7%EW�蟋�v��[һ��n�p��|Va�� ��ub��������Bg����q�ʐ�G�"K�����kxA�3�VXi����]��Z���Ff�B�����ȵ�
�Y��r�z��\�c�9���Epq�V��?qw�<x�n�$����>Y[�,��]������CED)nD���ܗ���dl�z���P{�q����\2�vcȞW�ߝ�?��#R�?!�N�v�͋C�>�H�'2`L%\���B�#JtKl)�B&��]���ճ�����'J�n����Q��hV�~�S{�pCU=� �E�5ۆ�<���E�UB
z`�ք/X[�5��qC����s�PtѰ!�#��'ۆ���Hx��V|P�9���Pّ�h	�́&3*Wf��雕jA�00�QIKq@�P���~d�?@��{��xK{��ȣ�$G�)��m|�66�7�d�� �vC�+���Rp~��+�=w�B��SS�_Ó[��N�7w8Kre?ʪ�C�e��!����`y;�����0��u{��vy
�H���)y��^����y%C�����z�P�y��6�V�kE���Ա9�Vo�v��/,���*�˅����~UJ�i�J�� ��3� z�؞���Sʒ�i�w���!��$�|�(L�羳&���������o��n�v����g��N<vZ�>��l�&����$��N����)(A��!��Q^ ���k�&����Ϋ옻R�.l� '��O$CL��|��p�zkP�$ ���]^7���hP(�������J�iw��k�l���.b�֖g�߬kK��T+�E:]T_���p�E�"&���@1�p?��V9�p*�p|�Cޭ]=d�I�6��'��\�>j��B�J��ч8�ڬ��9WQ�rB�[�˙��V\�u	�+m ��0ږ7�ԇK�t�I^.O�\
�,����b	&�15<h���}��K�)��
I~�NWtro@�gs�Zؚ�аs	�����D��`*��	F@M�"�_��mi�쯤	ٮ#S�t9�M�a�z�t]]���3\@[ P�j#�3csrp�٧�u�X@���T2�6pt�,X(��Rx��\���
Sw��.�s��������8��Ϣ*�+9aUUڕ�"1z!�a'߲]i���0}m5�+�]���r�P��>�"�"��E���#��s:��d$�G�F]_�֤ͧ� 991n�m/\sn���T��V�3�6�-2=��%=E,wkO��~�P�� ��$���GBSM<'�zy�`����b�|�p�@rٺ�TR�ܒeT�JM��ݐ�I���ut�%i ̺�2H��,�o?�f��#3��)��� ��Z�NU*O=t�.��zk�;�Z�p�O:W;ho^ȃf%PI���u��Ex@�D��++�V���u�k�(,�-���P�g5n��A��1��<N��0�����3l��a����17M�5K�24��Ɗ��r��F-|�3�+��1�
R��JPMK�r\Yߘt����E�o\�����x<��`�>5)����_#���ayk֍�#k�_�Y[:��z(�7�������i�*�7����⢺��k6#�G#���?��	�ԉ��{]wo��?w���@9�^Go�*���C23*x��Z]�Z�	x������_�MB/��4�-oq,�M�0�=_gpJ�>�mejא��5a<r�Q��aL^�����i��q��4+]��j�Y1����Lj۰����Zab�����:B�哮T94���4o�t�Qw��Ze�)��e���V6����l�Og��BR��w�,�^gA�p�p=I�rP)��^X�p��f��;�7+[Y�vh���-���Eʰ��F����A��w� �j`�)�#�U�LK�M@~]e�[,ɜ��ݮ�\�R��z1�`��S@(�l��I�o"���މ���w}�2��A��G�9��9�G@��c�|Jx�NWX;h�$P�˧����v���j�P	H�����r�Pp�E�c�Q�fZ�#�{y�!n:8å�l<���h�K��ە���k:��_P�&��j�7�1�K�����'�-O�A&��-�4¶ՙx��č2�����4f��]>#tj�݌�Ј{�x�j����g�����;(yoOۦ�4&'���⾪g��(d�؃Ȳ��}kVh���� %�k�b���bc�X���jw6JO��PT���NF��4Y�sƋ9�`��������k|�|�"lZk~\��f��r�������� �SM�7�{-��|��p��4>\�D�0M� ĥΚ�LqL��m���p*�����U��L9(@�c�lĤX�Rh�%S��H嘆ySh��P����p�?������ʝ����L�)W��gQJr$=y0�`���R���Y�ϲ�lS��;�.|�JS��8@���	˻*�dΕC�>^'F��"h@N,�����)Xvj$p�"k��A*ݥ�.�d	���=�2��ńR�?���⊠�0��d��:Ȏ�:�&�o�iа;��4�W��!��F܉����aP%�O<X����^�j[eA�Z�O#��z|\$�}Ob����$GZ{E�j/�5c�X�̓g|�Ç���U��)����Ȗ�o���$���+i�)�=��1x裘�}�I9����@N��N�l�L�7k.�7]���Y�ҳ^_%3��7%D�r 2�v��j=����~��l�|����X�� {�.��l}��ɉ��b�ￖ�GI��P�u��b㕋"&�8�9߽(óX1��a�ty��X�Z��@y�ehI����iDu��	<�K �@�I��#JѝC���&�f����5�_}��c<O�����Q�1T�2�����%�-<y�E�
˙�W  ��*�?�a��|{;M�s�]��V
�~�_�{0��HL��OE}]�Ca���x3�����:p9�0$Z��큭
��Me�	[��$�{B��2��G���0n�on��ѯ����V�]倭W�����^0���O1�ֱ�-�fǔ�i��"H��89��������>�+U�?.�9�s-?%ν=�!���:������~�X���๦6e�ƥ��z㚷&+ӱr}��߯��!V��C���3J���p.�R�+NcN�m���5Х��հ��G�/�?�����ͧ�~�Ŕ�c�Т�NӅrSAh��%]�^J�l7����[U�<ِ䖌<�������߻�Eۺ�G�7Y�W�GfUV����݋ 9�y�{N��/vB�q��M�2
�)����P��by`�sԖ�,8�e}����FH; ��3bn�{)�eK�-��h˻a�3.��tJ�����V�����M���bԟ�}�a}3Ƣ�Nwbą����i�m��s�ӬD>��r*�w-ba�!�7��N�X��cEW�@�]��$����m76Z���O?`1�%���Iq�Pee���̿�ϐ��"�����eE��t��muʢGc��I)��Ҋ1v�H������cV}��NZ���/���w5d)TՊm�ϔO���qV�[hZ�[6RAy�����w��AS����!+����J.�"i54Z��|�(�ir$_ي[�ܣ_�^蓐V>�$���ձ��%\H�����M���z#Sq P�/�k�D�4��5�'��3��<Bع��M����Q��
����	�5lT���n�zi�L' �����^�ؘ���;ˌS�����a��i�1z^]l(��~�������Z
�m,�3a�����# ��㭃���
���	pb��W0>.����T3�;L��h?��y���C5��{Vہ+~J*�@gn�� j}�Ŗ�L��{�B�ʱʮ��1�ƕOd�Et�S��2��悂�Τn�@V�J�l���Y������JA�3���|��7�I����u�����~'���LK�B��b��4qf�(��b�Xq�j�@�q�K|����GM��!��L�yN��]�:�#�R'gYk����,�^P�}�d��7}Ћ������wxKK#��cQ�z%�֨{1ʹ��rvӰD`�F��VX/u6ﺀ���Y����p��)��ޮwl=��8N���U���5
o���C��e�1��@���{ۄ��>���çS��]ȥ8Ԟ���ÖH��z�����h?��,[Q��j�n'0&�wY*���Vb��s�f��qL�sz�W�^�f-�n�DR�����~`���1��U=Z��A�%T:N��@y-�>�V��(]��
�9�d��W�!�3x�����x,h�y���f����L����?�=ft_!����p������1ñ�M:��)�]���%-�kg��=��b�>�vB|�]|2�3 Y@!9�Yj9\�z+ �kZ���L�QLl�?ܿa�F�d�u�R��m'PI�B�x�mV9K	3��;^�<Ө�0��, z�U���k��y��D����*���_ZH� ��$Iw\v��Z/7�6��,���D�P���m]�0�u�*�H�b�Re�j	
#���f��g���@��}sx��ذ��Q_,LPw$��v�Qyzk��M(�t"�O�AU&�w��]�Żbi�C&��1�*�V�	Be������o�bC��c��|�vkW_�j�"��P��@���A��g����{��{W;9(������P�j��8�j?��@�˙ �a㔌zdk�����e���gq8 W�`;��f�Qֶ/x�T�6���kuB>��%l��5me({�����=*����^5��9���w(��*D�D(2� ��佧����� u$U�؄��a4��*7kZ7��`@	6[��z̰��[�,�ᶝm`�X^�"���`��>OƆ
��~��׍� aF��� ��c�����;�H,>g���� פUD%��x�j&���ǭzͪzF7"�R��#�;>��;�32�m��Qq��69x��H4�L����ć̾/�<�4芏4�2|��:�SC�ۃak�5;�학!.	��N[i�	4���s��õ�=��d���+�}�/��,1��(�/
Q�[B)Ȉ)&��To�-��`ҕ����i/�d'�Ӱmx:/;[e�i�����6�7� ����}�ۤ��g�3l�l��X4���~"2��|	�~���<5�P��j��/¿L)�,�Y!�<���P%�u������H��x@�g��}��!Ͷ�S� ��NrA��[iFy@��$P�5��#y��qU�4�O�Ԁ�)a�	Hu�.5�9�l&�N���9�z!���`+����/�g����~��O�EڠO��7��64b�d2�(� j���G�Ǻu[H3kw�3���cOz��^�n�J-K�Z�<���CT�ܦ�_^9�{;OG�#[�=���5Lm�����)����|{��T�5/����(�����^3Vp��� �f�.�SL���$(�@r>�>+��9r7AO��T"�-%���[�Rv�k	�1����C�`g��(դk���i�r���ŷ阔#�1���Px�M7�m:����$�f;Vu&�������KO�1G�|��z#C�A�-釟�ɱqW��h�� 2��L�ȯ�Z�� �"f+�������p`�k�`&�^3j�˃=r�r#����ɦ�wPu�]��wR��v�)Ԧ�(�CC�6�2��d'����[~��?� G�M�lE"n�\2�"��Hf!��sz����3j���=��3&tr<3�e/��쫱	$բB�iG2Dza۾C���)C���`(s�����1�	���h�?���GE{�Б�-U��MMߐU=J����rb��q.���h���R��w,4���,	�r �x�!��49�ݔU�C	[�66X,}n�Ԉ��j�,oovf͋�پ7jǥ茅|{Q$S�z��8�k/4���U����58�"����:ҊP���w3e�L=��/�G��DM����w/S����:�!"��ji���ڰ��%��T�X��3d�w�G��v�Yd;� ?��2ȼһ[�ƀ�m��/Y���O �u�x��if)B���8h���\r E�����/0|Us�$�R�!�m�A�Do�]r�p�����&.�n�I�9*�l+��(�x"���b$ 2�In�E�K�\���[�q�0Uz_�=[�bs.0ɏ(8B�TC�;Ӳ��a{�a�0�ױ��0�=o����k�2bn!f���T�(Q�+���xi��v[o�s	<E��1|�f�9�g�,�"(݇2�#l��٪b�Ԛ��I;��Q���:3g�f��?��}K�J5[�=�[��9
>U��<��{G��G�8��._M��a��㍯�7��~~���-T�<!1�齄���u���GXY��������&M����%���Fhۘ���B��O:��㻡7%��:-�b$�|Cʅ���o��ԎƕY_'��
���=0�v���]KBoMӍ!Ӭ92Xl���D�����8�:�A�g��)�NC���\����ww��zQL!�US��'G���ҝ�ֻ��2a�'����s0���2�[���L@6��h�	�N>�Ռ�����M�խ�Y=\#� ��R��6@i:��V�ݘ󏾊A���#��F�?{�keY�s�=�j�`u���{n�C`��F��3���>�P4�B���tgm�< �U�R�ǅ��g
7���h[3�NX��'v9X)��wc����T�5Z$���zש:Qҙl-S��cEҪ�נ)��J�[�ʕ/b��;n�O
i�t���;����.#C0Ґl����'ll콘"��i�C(�i��{q�:���C�@�x*�稖6	��]�)�BU*�s7A+�s+�������kX1�}逼�� j��+=a��2�h(D��#��v��_��q����0	ګU�4�z���?x섮��qz��@�Ļ���V4 d�:,�V�wBA�6�0-��N����ù�%$����T��w��v��*���r��{����M�卛�{i��4 �r����jwg�耏�5 )g�$��t�rf�X��7�Q%�y�L-|g��Kob�hYF�������*G��Y5tȓ�!v�0���Y���!S�7��y�H�a���H^N��Ҕ�����R�6���&8�Mv��MZL�>"�<�q�e���+�ѣ�E}�R�`3��^b�y�R�j4E�^}�9��6Tf�T�1B�	��9t�#f��\�p�
�
"�����ta�ō���7�פ)�u���I�qi1���P-�ޣضdLJ�a�Њ�+v����f�F]p��[�gFkO�۴Fa+=N�,e!ϟԈ�!=mL/��-yؒ���9��#A9��sm���z<�!�o�&D���45}��"^S��鏖"��lߓ���p��q�8V0pP��FP�	Df���4k���I����?��b�M����aҲ8�;y���]Д�~pg��S���G���%秾���	d˾}n�!�R�p��^A�J˅2��O� c�3�\��j,vVK·��ylnꇋ�[l#�rZ��G��_+3�=��;.Fx60H��ݹ��t�-sh�
�,���Y�P��n�^�ZR�V�N�Cl4������&4� �0�s���{0_r1p:	�C�[6Q+.� �Rcv��V&�Å���08D{$��C�&<O?��ePUW� zO!c8?��$N&��TW��A�� �0��q�
G0��x��~����R�sQާ)�׼��� ���~���=�5[Uۥ�{���YeͨL���$�$y݄�k��Єt�M��j�Σ5���}"�.�xJ�����޷)��(���4{� ��/���Q�z`(<���$�:o�-��Q��S5d�R����c�ZqE�=�a:>m��Wnv�#Q-��٩�8T�4�@)��u:���Vj��t"�n��4�J�)��`��xq���<H�	��p�ui0�D���D�2�Ptb�zA<��#��$��K���,Z>1t�S���h�L�f�i=pW�rl�麟��x��I~;)OuM��0T��-m)�i��n�9iU�X�f��ύ0A1px�Q#�v��Y�hbS�cr�W�{�b�;ǉ1��uӕ��_��ty��u�
�&�M1�l���� =q�L4ลؿ�1�ݟ��U�������ɨ�\�O��$`�ʱ�4]У�xU�Rj�;^�.p�_��]6��Ʊ��_���Z>��`0 �?"�ӽ��./
��	��K�@��� %�w��Zxl�\e�;���m"��+��qL2A�2r�*��5HMk��D^5;=J{x�ZrDʧ��k�n˯"���u����.g�i}���ML�}N������|�������?t��	A�1��#���� [V^Aa��7t$zdPO�兡�ؚ���� OWK�uv�V�n��"6t���O����4|K�X�bB�� r��h�h7�&6�Mn>�Q���aS��HY�t)��%��| �#A��z�ڲ �lA )��\�\�e��NYΗGlBӝ�������Ε����כk�W�� ��8����Ō�t���W�)<����S�a��'4��K_����5�_͞�2�o�"���b١�ђj�迣P��/̟�sb�(����'�Ԓ5�Q�R��EӠ+ȭ`A�B���1�2S�fB#�-�@�H���X���+��u�b�Q8��_W���I�
u�mN钾D0�巧����)���8�FQ�B���M��g�
��L�zG�1&��c��^��3��o�U�Y��>>�:D��+~(n���[�N�	_����}Y�� ���]���_��i=I�A�i�l<^�k��
)����>G-$6n7��yށ�ԣko2��">_�����H^��q��\����"��T$F��~)?�=G^W�P�[�������0pj �P����
L(�aH��?sE)����ԅ>�Lû�އ]ci����P�ȉu鎗U&��F*|[���&	�\�C��'����[�P����rI�3��M��R�*$�L�BA	�M����ja��3a`[�~�-�~�D,��i%�nr�	5�n��ˠ���$�|ܺ��߆���x BhH�!!�5�1�XG��0vDS�ў1�|i�kģ�������?NGD��4�@��K+��p�[)-�Y���#"
�1�����7x�)��i̪��p�OYB�Lψm{��f�}9Gy���X��_Nu�%Be��毳���>::r ���+1%b���ۊ����\��;�����E������-E��2JjO�۹�m�f����+�.�.�B0d0��;F*�Ε���T�n� cːya��Gh�_�!��[�������1\9yBV����\�4��/d1��o��;Ӎ�hoD�\�ݩA��'﩮�5�T�J���҇�!�D,X�$���B؉y��osT�C����qm��v�j59�3Q،����K�@O��v.�p��<�������Yh�BV
)��������� B(�㎏xw_E��z>�jE�Ho�aQ�8�H���� s�z?�7����{ƭ���	���ҿA��IN�G	hh�ӈ���9r�e��\U��6 �R�y��Fp�К��q.�W�Z�qK����Xy�]%9��ڽ�g��a�̖�����ө6_�T�'�&Z ��AzÍ��,W�$��Zg	��X���F��=����w�'!�����,m�4dJ4�	{dT�����a��Wn��������M9Y���}��H�\O�X�(I�΀�b�\�~~���*P����a��C��r
=B�:@�R|33y ]���܎��ǥ�}P���py֌[�mj�����u��6�@mw�z�׃՞���(��R��U�d���?+B* �?�k�1����N����r	��� n�:��OK�l��S� ����B^nӦ�l��E{�D�����{#h�5
)E9��T�d)�������;ǲ��!(Lۊp5CA����ݎC���G*k��4���(��BC��0��]6���x2b�&+v݁,i�+�]��k%n0j��%{z�@έ���Ǹ 5t���N �@h�
�Ԯj��c����:�A}
�n0,�t���������w߷$����(s�Ĳ�c���Rh���V6!+mNV�	��}�fJi�]��G�A������%��EAO��@�����eT�B_@̴y&߳����+z�����i��t�JS��̕0��~L��z��@�=����JH�;� v��,��� [�8�ඎ������
q;�N<���E����-�)6�@IiK�w�:��U6��\��kµ���X&̘z!I�Q��1F|��E(��v�f�C�-��))�h�� �6.a��i���?P�չ������Ս�y�FC�ݾ}O���
��.�i%a%�zH����,/��a�_�8{~溕�R��y��f,�j��6%���xp�=�y"�0�U�� b��5E#���s�B7K�O��f���� {��C?��ɑ?���z����UP*8�d�@��UbƵB���U�DF��5��ɋ���I0����3V4Ǥ�N�A��dϒ�p��AZ'ĢM�4����Y|LV]q��e�W<��<�q��j��)����?2S6Q�6�K���8+݉����,�!dwvO>���j�wB����׶m;��6�T,���k6qu�!U�r�nP�ymb+��,6A�zH	1�wU��BX�����pV)�oLn�	莠]B�&iLס�}�MY��{dhӃ�ϴg����:6�>��H�8�1�G$��Tv^��'�tY�<A:�ޓ��%^��;~�o0�E��ȡN��3�=�S$�V�GUR�����3k����}%v٩��*�7��W��!F�,�5�Ü����q�	ǿL��2���h��m�Z�I�Ov��]��Ӭ-���Ɍ�b��m �F��3�C�����6�z*�1e7����g�'NO�u������+�E��0�v|��1������z�@d�a��}D��P��0-%�@!�]W�k����r�U���|���̎�ʊPxj��7-Z�9�{�K=n���Gq���ͼ����C���ʜ�Vϔ�	iC����_3K�$YT��hp�� RFZE�&�A�\:��<�`Fi@ya�9G�`_��b}<������-z'^�����'�h*q�E��Is�n?���S����z�k��Z�?�ܸɐ���b���R|6��K���@G��	Ό!	:1Տl�:����!���$�G��3x����Ҹ�?�g�u|v>u���nV
����			Q�}��H؃��oGJ��[�����J��*�|���\p���\�j#���wi�Pg}�kWh�I�(A4,����0��C}D�%��h)����ל�H�Mn���������X�^�8��?Q6�p��>9�_B�+y��&�\��b� A���j�؏f����}���f������^�!-K7~u�b��lB���\�\�%m�8%�L>&�NdF[���ZSb#�#�s�s%s�� ��d����1H����{4���Q�T���#ӝ���;�KBڻ10>�6����2oS�f1��(�����"Ti���Hq���B
�#/�"�1F��Qb�aNz�	�(������p�Q�}�/�ҿ�����S�Ŭ�'���t�<��f�D�A�O5ݜR�Lv��nA$�v��>n&�ѣ���¸x��'� ����v;��%�"����m�����i�aUe}BPRE�8$��p���c'�nHjL� �%�UX�H>Aڞ�o�σU~�
p_S��EBT2O���K*<���W�LJi}�垶���-n�T������U�����ǣw|�Ǵ�J��ǣ�T�_�i���d����5��Xg0��M9�S1|ֿ~��9�;�7���<�X(�u��!���6�[�TA��_zF��T�P$aQ��
�[���>ɖIm�S��ZنF[��8}��~����( c<��^ƿZZ��u96����4�7�K7���{!(`Չ���� ��e���!�=�ܽp����;W�59�ad)f���؞�V�K�VC��*�w���iK��JG�^����s�߽D�n'�#�JwL��_��-Cm]e�~w�x=�+�#���3����c��X��V=�������ف'S3����'���Z�/��w#X��)���ߐ�J�@�]��q��F<�VT�Z��n�Zz�}[�4�@�>�N�!�.��pa�G	F(ф<�(W�������j��BO�fϩP�MBO'��Lw4j}7i�A�@axlɺ�WޓġT��
��K���ľ^L�����)ߢ���IF�Yb>�!@�&��S�ip��O�	��aLN�����I=��Yxr�ѽ���pcQV`��8���13K��5�,�{'j�
���q�X�v^h��s�#�>Z��m �C�O��Z�.;��|!��eU��F5[&�QɌJ(J�Z�[;���d+���~w�j���ۖ4>c"������Y�j�;�����Z��X�~U�e|��C�s�:F;�r��x1�"��0蜊o@�f?Y*�_��N\v��T�]T^Q)9�1[y`qn������Q b'����_�����R�N[3IK�"�x�:UTQ��ir�o�.(	�ӂ�APO��z���Df��N��<[|XNnp6�ܘ���Y��ʯ��{,'������f�:Oo��o�޼yڡ�V5�\��Gԅ|Gٹ���Ά@؍��*k�����Z�5�Id#���#o\ZB{���!�1�d?��b���G��>���ew�͈D��0��ł�aeR^ˢ�s�L��]���Z8��~y���3�5/\�#3U�3���e5q�g����mA� !ə��P������$D���;c�`�9�?��E����I�؃�o$ì�<L�O�g}JBW�~/�O'�<c�	��_�<?oZa�4m[��2밋9?���� i �Ϲ*�	5^�d_G�wU'�{
>�j?������;�*���,��$���]������+`Z���:m��*�+�n���@�%�&�e.�?#������$�n��j�{���9�w̃U���5��� �m)b�X�4�m鋬��;�;\�q�^j5_��8�nT��jb>Z�עP&�,tӣ�S�%7.�.t��
p����#� ��(����Un��^u �ڠR��MO����`�ke���_<)%o?$���N�K�"��#�^�����vt��ó@_�{�r�fy;���^w�eU����'���Ma^���B��ڛ/�pT;��J5G�s*�5�(��H�����&]�`��x�m��!����FE<V�B��x�S�5��S����s+2s������i�ݢ��Z��Θ\�$���1OoS�����q���fI&R�Z�r�W���ml��E��^S�������&��Z�*�1�\)+X�Ƞyz̓��5:�#���#S�w�����
�x����~��ia����x�S2#����M?�ˊ��t\%d����p��5z�.������;��t��O��?x_�K���Z�Y�?��@&���>*��PV����F�j+�ֻﳶ+�p|�-0�]���z�M� #��F�<�r���=D�m�t���-v<	�/Q�xw�*���r=*�-�� �H�Y���b�@�Ek�q�b8q*�ˡ���V�?��H 4��)W�����֓��spn���<���#�ɔ���]!C��}�I�`w3��j�>
��������٫J�8HS�m�dy��a�+�r;>��*��[�QC1x`z^6	m�|���D{��:(YBdy��Dw+3�h'�M@j��W�~^� % ���GB	�/Z=ӾC�sӏ�Luф�l=o����=�{?�0,ź��D��ei7�DY�;�Zѽ֗~TS���Mý۲^<�y�y)�{�NtK��lC�<�1���=Bk`\��w$.)Z���66/�Z�"ψ��
��a��N���y��`K4���8�3�������0C���ɠf̤s��F�����`@��g%�ؽ�`2�$�Zgr�7�D���d˖0d�����g�Ln�f�c��E(�SBNFr���D���l鯴��Ӣ�<����ڨ�_��0�B�&<�f��G*�aG�g��9vن��G�X��%�����ɀ^�m��U߸�Z�P�I�P�#a\
��P�#,�!Fe��%��t�� �v�m��U�-�2���e�����g�(Dd� �?���KDԪ���0O�����2���i�51��� ���'�Ԇor--�2��z{��[j=��Vߊa(͛��bl^x��gq�r;W����n��G�ȍ�|��r\����SY�zH��x���[��7C�&��
Ѿ��P7ǉ��]�	�CwSDF��#�Ha�`��1�k�|R�(�Qw���r���ɻ�ե�< m�nY���6gXZ��ѧ�Fz!��J-T`�U7��UӂtF�YRtL�����>�60��ٴܲ�L%�랞N�J0�� �,�rϬ��nO�����6@�ڋԞ�૶\�0Cxآ���Wj�?�Ow�z�L(P�hV8'��U_�1����%h	އ*r�ˈ$�&�E�>q|�����
TUf��i�;o���pp�+s���;��� EڙW�l[�2���3�T[��*~C�ܐ�~d'Y�${J�[�2�w"|_��l�?�7�{���ÕA�q�w+a�e2Kd�0@L��9$hD� ;��r����;p�{D�9�z���6t=��]����<{�8e�[��H���o���9���i��ҩ/G�T��'<#��q��N�p}5��.� �6T�~~	�l����Ng��qh����8��07�ςϯ|��S��o�F�w��ں���M7����8:�L��t;�X�!���>]zj/�Q��S�E�q#����>bQ�Ժ,l�ޭ%@h�m!�M�'�f�I<r�	�@�>���f�Ӌ��+�����Rֶ�%)T�A΁��a{��H�����	�/�E���!��m �O6��o�|��`Gy@�HEu9�e��� L9p�<?.���>}��2gm�}$36=x��i��y�[7��D?ld�\���!2���#g�2J����N(VH�#��^��
���I$���Y&!��{Ȓj$�x����G��pyy|��)�<�m���WK�x�����w�(�NӬ�Ґ�*����ޠ��_�=L2K$!�m�#��C�пԤ
��%���V���PZ,�##��=:ە$!|�h��}w��D�Rn��~F#�A���-���2���#��P�����{쏡$��8�j�D.{c9��y������*p���|.���I����/�ṌMR�������wp&.wi3���Ϡ�n��Y�v�M1R2�LW���!�L]��ك����Iq"q��3L�
|�D���p��j>���*@��oUy�H<�C��.ĳ�LK����j�A|&� XU�!)p��>�gC�5����b}�R���q�]2]y�Gth�4J�j}���+�/o���C����zҩ�S|l�t�>H�'9�.e����^zI@��&�u��Z���m����ӌ�j�W7�} �hP���D�gL���8r w�^�	71^�e����6��/
���fV;*�Ga<�<3	�o1C��M�P]9q�A�����M�l�H�|��:@C�E�]m��G���AC�r����%"�R���?����Q|D�ij0.�!7�w��JP��u���cǲUJk:$Ti\�%�W��p��{�H�!�Ge���uR�L�R'�3jd�⇷�'T�WV��㥆��R���;��h<�L[�qG��=��B��:�n���#��n\v�Ϻ�
o�J�o���g[v����c��l���>!���'gz$h[��8����]��^N����	��_Fiv����䯆Ȕ-"���jI��eMM�kO����E��[ v��<��L|)o�@� �/+,@��5���%�"���+G��s�N��%G�g���Ѐ{;Εh�}m� ) Mc!B�.�*�[��=��mJ ��#�u�[�8�c8�k�=���0o�s���*7��J����Mf���,�z���H�"�x	n�?w��UKO� @}��Ԃ���1j��U�J�nۓ�&��.����ϥњN�]���0����r��*E���:4�:{�`�_p�;�8�����DEe{(��cu�ٕ�st�r��E�'����>O�m�̶�76��Prpx�E^<m���1޷�X�m��R�z��:Ŗ��0j;�g�_�7�>��ܳ]�FÁ��dU��Xv��x0�LC���-� \����v��[N���2-�=���A!W�n�$�D��yB���o��!f���K�\0m��[B�sj�3�b��^������X8u�M�;|d&Y�<�u�y쒢��f"��$����<ȳ����QJ>YD��f4p��Vp���
^Xk$��P���z�_Br=����#fAǪg�u��B���
cs���Yz�!��l�l��-#/)�4�ڌc,����a�dHWB<bp��O �K�8�E�dH�;�� �W���� ѹ���̫ITF����}��b��U1Ꝓ�1�v�������P�[�S���p�4]@Z��C���q�}��Б�o+��I`"J���X��M���&�ՏAY�[ݰJ�4?N��㺀�Ħ(c��e;���*PLm����m���`�uoW\҈Ktd�i�/_�����R�K٢њnA���k�?��Q�����ƪt̄D�o�&��OXMre�G^p�R�
�8�ݚ�iWQ��M�cd+B?�� #p)��k�N�4\� ��&B�n��(.[���H�̯�$��s��o�Su$[�zk�]���M�=V}��K�P�z���\��m�&>�n{�b@����o�&|���Ҙ//�*6p�;����n���O͌�y��Ӕ�w`2��}�,�Z�`�Gd�P.Ϛ@�H���Bp"�0�a;1�7� Z�e�Q���\�ݑ�d=����	c�������ѥWT����B�����s��6����+'ي+J�LUm-�F�>PJl�]�4�� �L�*.�#���y�ܯ-�~G_-VC��;���K@��L�{��ج���h�T5eN� Wt1`�������m*9��aod�j��5����-n]�:~�����O���^��~C@b�����T���P�<H:h[�^�|1V/ZvP�+��چ���z�ʗ[ْ9��R6��ҫɪv��0|R��@}~���J��u����(�R�I���&��s����������-����oӵ	��USB�
J���6�IVf���!�(�X���� <��$���9����h7��e��KP�[PR������-@K�_>��c����j�>K"��2�����������~������������ٜy�}&�sPĜj�������Ү��T����;��Fx� �]I�b� \=b	��u���+Z��@�_.��%�=���>k�������GHՄE��ʹ�<����%��a �p�AX��J�zKu���茉V���"'-Ħ�'7��Fh�]3�B�q��lÂ!�P�
K(�Kj�P�5k�ޑpaD�����W.��j�1n-߷g$���z�3�0�ZY��r�c>N#�h*`�<�T���#��1J��Ǆ��s���oNZfLG>t�ꥐő��7�F�XL^Մ��rC�d��Y�nP�x�,��������FJqQ+��c��sh��KMf���#�/��tÛ���qqO�I��?��Q�Ε#���H���P��[xK�κ98���u[���Cs��ݩp�"|�����I�͹ey��T�'�k-��W��O�h_Z�=A=~�5S��7�.��3.�Y�{�^�훡�X+ȋ��oӷ�~�k���Y1mN;��P������Z��I�/���Ƞ����;;V4֎���@q�jx��/�n_�Ɍ콭��L]F��c����9.���=#� ��QӂZ�E�"s%�?�`��4�H"��| �l��H�Ak�=׶�Ξ������ȩ�5���!1��^�O�C|4�X���ȇ�6W��Ԗ�'�����H6.���}l�k~`NG�u�B�`&�x�=ٔŮ6U�^3Xt�����y׋s����L�$�2�j�D쮷��؝��h�e �Z�jթQd�`����N�e��xr��F(AnD$�R�M^e���H�-}����� m�ǝE6�(�=F�`@�r�w�|ۗ�7bW-��*C=I#UO�3�6�W�B+Hb�LU#��9S��Ux�W�6��Z����Ԁ�q������ֽ4���x���_N�?~�"I�7�Y&X+��?��Uf(���ze��'-����	Bf��(5�א��v���]�^�ސD���6�0A[�z$'䛣N��c��'���:�D��+�8%=�ug����e-�����8�����\C���C$�Ⱦdt��-�1[���G��ʨW1Y�Ͷ#U8��"1��l~�|fq`K�rWܔ��QA�Wf�v^Jw)L�8����֭;�B��Չs��@G�gtxّ~n�a�M�$�G�[^�����O�QT@c���7�%��5���X}��at��&���I ��Z.>Z�"�m0h1��<yН�fߡ�r��7z7����MH�2wJ����x8D�Q'�5�\��E��v��!��]�O2,Gk�K�XGt6Y�,�-3'�������:ݍ�UiZ�z����n�u�"����꾅�,!l%�����Or#��t*�׭��J����_7��\�\��Բ�_�KO�-����	�O_+m/��q�x1�pL��OG,��Ү Na�K��ڇ٬�X�8}?�a���ٙ�7-�����p���7���hI5r�m�O���wjV��$KIo<�m��3�	�9(]�k=�᨟�� T�b�Y}�f[�U����G��QV:07�2�Y�������V�9BM\�3�ж�1%�ꩱ���.�9��-
]R� �B��A-�w��� �'d�������9�i�U���ϴ� �j�5�����Ԓ�U��	�q�<����1C�su��2�=��ۋF���c��م<\KI��E� Lgޖ5q[�,_U��9d�1D��Lw�6�>��ʩe��̹�X˻�O�����Q,UA�jJSg�h��zDd�, U��*p+f-�A�)���N�ښz:ܩ��ܙ� ��CC~4��ɜ~�~S�^d=�%�r����cQ�Y�c2B�h{�>�[v�K�lh���;�m�!l���#Ah�4���T>��R�_�h0���&U���u�9�q4����Bͧ3 ��5�/�U�>t�ҥ-?���	y{�� �Y��5�lt�E�,���{�+X����m����EV��%젦e'?tK��W6�GO�)�uZ<g(���U�P�ak����,0��Mjl��#<��`�r��j`�0���"��Ax񕒅����K��U�lWS���ӣ)��퐆��M��R�{�tڅ�]R��bщk��_��!�|����R?�NX�|��{I�6pb2N��h��Լm��L�s@�=����tG���Ec�I:��8�L�y�󱾁��2�@�O�2�^-Is��,�gէ�wJ��'B�P�u�?mG�[�"7F�7	���N����;���٣}�k����jx���BH7h"Xp�C�c]3�G��`w��iW���V��
�z�B��1��C��[(,�y����9��7�7���C�}�E���߉�_44�
�Y���.�4xD�������g8�'t@�6���/L�ɓ�E�1���=(ҹp�q��*Ss���q���E����i@<�S��`>ϼ���F��{�|g�/ܺ�f�����j_(U&G���o����9��<���~��o0�x�8S)����"�E.1q���!䶡=N^���S���e�����ш���ƨ�g��|��{��Xmk�1�dp%���j��B������8��[)���i�r���! �s	���[�%J���Pp�-�x��Ө�l���mð���ah��;1&�@�7c�l��������E��e��>�H�d�Oڙo���S@1��ՍѦ[�M��%+LB
+/�|?*�|�$7�7Q�  �@p��b=�p(�0����Y"��*����O��MQAFx�/�d	�ą�,�#���.�-;�b��3�'����kK��*�"ai@L���*9���<#k#(W�YH�w�����Ր�ϱ�+d�.���N�b��U�;Gt��.�,��*"�V�r��x�73��er宝`P|&@�>V�G�Q�_% ��N~�4�/�y���8SQ�gHHߝ��6x�k�.iRg	P��i�g�)���z�9�(�\զOk�	`�H,�N�ĈU֪_�UP�\��XiɗF�\��'�V����^����#w�s�Lcp`g���J72!ME�׏��2�PG���6��/�E	c*�F��M�$�ڻ�t[�kN�1)�6�1�c.R�ѡ�xa#�m�1�pC�(K��ךuZ��Fs(�.a�~�������7LwS�T��Oa���/Q����q�*��ň�F<�����0��1�(G�$��F~g��L�����!��6�FI���cd�1E(^#֒nI���`��.lqC����#�-'s�����/軑�����c��L<,#�q�
��cwR��3S�?m����`I��M��]#�����eෙ�ok�����Ӷ�כ�:.��?�(*±�`JÛ�1�C���Tf����dޓh3��PL��
ӳ�ņ�c	�ncĂ��f%q(�N���р�P�ʽӂ'��+���p�`H{so��=���*m-F�X��C)��"i#�r^'��R*�/�y|��-fI��WK
�8�O��}Ɵ���^U�V^S��qQ�^�S�&}�����G�;�tU�)�=2v"?Ź�d�(m��b���/>��G9K� ,�1�ѩ �(q����봕RK�}��	Cu׭}��%�;H�4�r�Jh��wd�������b�M��9�Ҙ���v&d�� ,���kX�9Ht�ˆy�2lv�ձ���>7�G'ө��4�A�>|M=Aa�fX�ެM Rov,Dzf�YZ��CFx��Y��S���t���A��Ӹ�]�]"Ϗ~�8�:��^.EW�N�	?{^���L�,%g@������y�u�Wgz8@�� �5�7�\�:,�G���iv�W�M�Nur~�2 ��80��_Q>�!�^�Ň�C����.O���
�S�S�j��T�i�,�h��!�\u#7��I�QW�L{��vvsB�0&��ˠ�h�'=�Fy�n;��K����v��\��k�sC���C�Οp����"��U�y�s4EqD?���l��sb��:�W���vG��^�y�����Ql���]���d_ק6��Z���F٦�Z�Y�L�E�A��������.~Q�x��P���O������kIvt"IR�x�qA	��@Y7�J���tq��OUz��[Mnq����1L{Մ}>�,4���X�䲳n��B;�x�>�΄��Ha��<G�m�{*�����z_ē��ml���!Ԝ��1gk�O�:���� ������g�+����:�37���g�y���zuA=�a� F���SHM�Ll����{G�v�{u�E�5���а�:t,�W;Ie���������moY���-B�����g+�"f��Vl-���JH�!� �O]H�lwٱ��eC"AU�Z��)@%qo7ə�JQ���Gu�=�tYlD��(/�~�?�h��7c�� �K ����I�tB��̑�F��v�_B�Kys���}�[�o�~��&��d�4S�B`Z�]�#[��4e�[y.u�=�cJ�"��x�Nb�Ŀ1�e[)�M�l �s�	�'6�N��Y&��c<d݃�Ë>�>��G�K�;��"�Qൗ*�����7vs^"~:�|��Lp�4����.��������[fD^��{���Hz]�_(T<�8�����'������c�:��6P~�ſ��Z�}�F����Z����v�y�oZn��o�h�{W{��£�S�-aM�u��܌�b���}�;��Y �lB��ϓ�n\.�+-J�s�p
�Ջ@FB7s�D���3)$"u0M��h
U��L��S��U�tG�걽�{�c�|��`Q�
�Io�0I�خ�{f�x�5���n����Ԟ�����SȊb������-��y4�{��:.���is�&n\�[�R��p<�k�cf/���g��ͺhu}�n��6Ql�U ]�f/X
�孬%�1Y�p޷]�_`Y�� ;�Ͽ%�xqL��s��lsFp�-��A� ��{b,7$��^��HY��<��ݖ�x�d~yj�Ǹ!-���F�&�qLN��:���J/q�9[#%�N^+�%Mߥ��|����Q��~������u<���x0�>n�y�Ձ�\�`�.i�J8��\S�E
mtK-r�V���)��J�΋�[ȅ�A�j�
2��.Q�^r��8 (^ƴZ8"U�n��RZ�WK�O�!�	�5�\����@�'t�:���>��=��];�ɏ������;�̿�\�2ə4��1�@n3>R"�[�����f������~��!��� %�Hڲ�r��,�R�%����<�q� z��Lf��0+��,_S��;��u�(F��W`�S�w���7}tJ���?�c��ՒѥP�9���.�z�;f
Bۺ&+��Ȝp3�D��!R�m@�BGr����B�#��� ��Ah[ѕ*])R��g$hY�))lE
�Kڔ&��&�PR'�����/�%�LŵMN�����S=Ҏr�]�l�/|�+�A>�G���Uf���O ����ޮ̽'�f�u�>�_`�[� �Kt�U�ߒ!*l��ު�fG������6?�RR�'�|"�h��'�oA5�1C�d}�I�rJW^sT������&,q��`�!Of/�n��u^��[&�6`QΘ�k�!`��m�<1�a;ZY6Pו��&��\��R��G1ȷ۟ ��񚷅 o_��&W^�
g5�P!I)��'�?[�ai�ٟP8�p[��H��4r�J�% �&�w�=�߆D��6�D���������VG� �� k�����Y�m'���&���N/����%C5��l��=ҝNV0Y���]��ї�~� l�sN��{o\��ĥ���C�<��
8�W���y[W�9�Z�\r�p�;/M-�q����+�.%��:$�����|!u��.�Z)�#h����_J��~FN��v��d��C,�G��e®�����,_#U`�:罢H����h��ϰ�	������JD�3z�����t)�Y�lF1	Y����������^�6�����_|0�~�&�6�t��O~�m�фD�_�� ސ���K��5a@��gL�xT�}m�(�Pd�-�Њ�7��ʅ#�Ou9{O��YK�r������̡��JB�#w��"�7����b���vzqF� ��B3և]��>پ���
H����t���_iJBiOKR���r>8�,�v�����B��>��ֵf�~�;� �'"	�N���ٱu�G�.�)�]}�?/�?Q���H�5q�2y�����E�v�޶�x�=_��\=�v[��M�u��Yޚ2��my�[�>����ev��!�'V�������m�'���L�~<ƣ�۞�>���Ǎk�85�����e��E�N�XH-��|��A������/��ѽ1���M���r�.K?�?�pJC��t�M�w�)'7�u[?�;����ߡ�(�����:����:��T���c�� �9�a����X�8f�����{��XDmҒ�M�d� 2���5v�M����̩�m|-�7���'�T#�+���D��J��s�1��G����r$o���X��0���O7i�x�z�P �s��u������ľ���uٲ�Y'�xj�w9K��d����,7l�%�3�\b�:��p�yx�Vz>E�&��ǶnMu�X^��(�~�"P#
4�x#(݌"��@V����7���z��� ��r�����S'��5��t(�]D���/Kŝp?����xh�.1M�z!�&�����FȡF6��\/���=�Jk�68��)���aF�����ՓY)�K7gUń�P�q0���f��������L̖ڄA)a55�o0�]S:�5RQ��:���2�!a����X2�WR5�z�������7�f������ְ��D�M5��=��xw2���$�������c�'Y�R��ܭ�tj�^�B������{	B\�W�TMF�^������ڃH��o��P�q�V#fM7� ����dt� o4��J�t�W��f6��)�+��Lf���?Ĳ)�^`=KV�9O���u&�a����i~P�!�
��*K����u�L�c����cu+�RI�qU������fE�F`�Py����\@Ck��쿆���������q���"9�4L榑���d�!�*���ʭEH#�6D��+F�b�T��6��4�,eՖ���~A/�)�!�:a(_Ү��yc�Z8��Zsw�����%zLb�"fv:Н+���%x�fU �� ��#Dl`��.��¼�����cl��p��i�5�f��␬ ��s|_�(��{h6��*O8i�C��}������t�0c�aZ�o��R�[PgUY硛jÜY��K�`�ڀn��L>�B~�%�����n$[q1A����f�1�&�K*�WXB}��9}����|�2%K�6�ˀ�ؕ[TI�:��1e��92��ΖM~Ȁ�Q�h�ٓ���CڴD�f{7	���_}*�	ʭ73Xb
C��c�Wҟ�c�9�6�(���/ �2�M	���	M�R'�b4���/�E�ՅZ�Ek�F`��R�\�SGs2z���3w�8��4eH!��O�`��8lF�>���ə�t���m[˕w��5��	����ZC��XI�$w��fx�h��`�>�U��y@-�)�^�VY,A���'�#9eyX��P-�u�@C��l�᪜F�pDsYU�D��y?�}�^f�2�ʯ��P R~�@u
�(>g�	� !�6?�0 xTO~]+w��}a���N=�ꖍ<y;�����\E��zm���0R���ml�����w�߾w�++ �G�킩L0U�~v�!n�%NT�MrV���	m�-Y��7�6v�q���ꍺ�UӼ�[��4�!�ʢ�$�!Gcwo8�N�0r^��n�:������%K���e�t'="��
�N	 ��~ٷ�-Kl]�0�M���ixZ��kc ��ix���2��K�WK44�γ��'� ��m5P؞eL�V'�q���:��vU?�\�\V�.M(��@�������CA��m��+\0I����R&�svWx8O%9�|�Ί�Ft�$ߨ�f�'&�U(��W��>��4���h�夳�E�F:t{l��yz���S�[)GF�}(�*w6B d�1�Y��_�y�c������Y�R(��m�(�۰��S�m�f��ܶo+��e�f�-b	4Н��(kBk:��H�+g�k/uI��G�=3J�Vm��Ѣ~���k4���Ε� �La��j}�yb>�œ��O��Q��C]x�j��M���������2�U��}�"Q���1ۣ5�-ʨY����0��f����D��F�%�� � 4�;��U|�����@�y�^�A�4�k3���U��] V��
皻^|���%ȯv�ǝ�{�Q�!���F���c�q���l�%�2�I6��p]-���G�����ʅI�Cν.3�T��Ƈ�e�txQ�b��Έ�Я��~K�'x�� ,�[��w�
R��:+Α����ENlUw֚E��^��!܀O����]:����ԫ[͘�+-�q+j��g�>j����r�g�������F'^�y�v����k�S@6"A�/���_2c�xo���8㏯(��>YD�����!|�������s�aϜ���U"b<$���f� Jӽ@cU�E#��Ip���Z;�\f�;�Ը���k���{�����.8�{��j ��P��м�9=���;���UB��u~U�5,O����l��x}���z���?�9�U?�L��O��KW�B�j�E1_�G�*B:65���I��E@_3و��,�^D�F��5!)�w�U����kU�1��Y�l�6?��� k'm+��e1�|���U18�C�p��)Y�#�fQ��h��|�����~�%V,҅C�hX�7˘�↶������t5A9�l���	�P�:+�+�2�~*i9��u�q\�g1l�\� ٽq����\�P'`���_�W��Հ�@���Tdg~��j��m1߂�:��'�#=w�4���3�u{oZ�HK��ӽ�.�z��D�T�vs4i��6�v���u�3��%���~��*h�2�k��Iq+��r�����G�ao/(�u��AJ���߶C���E�Z�1WL9�	e�V�C��v�eG(er"U>�Q��4�F���;��m�'ΆD*�+B(H�I`���"�fhH��5+Lݯ�'�Ú���Q���ұ]�������ލ4��C/�m����S0��u�3ga�$��B�m�! ��/���h��C$�lj�M��`H�V�.a��N���1m���??EB��)0�L���/@"a�](��Ѥ�q->	��l�V)���2~�[��	�/lօ���l�-�㇒�>�׋�u�e3�
��}쬄�7.�ƺ2���5p�
|�ji���}�sA��գ�GQbC����zг�d������"&�E���6�����Vj�k�����T��L�x�e2������mi�@v��H^c�R�K\��6�9�\B��_*%��U雦Ɗ!���aH��S{���^�\�O����EC��N�z�̨X0�S`�4$��?*�*%����ԉ��M�_�ü�=�䥫�AE�9!A�@(R������i�m�+.X�y�`�Gk��>�Q/��Gк��Q��	�D��Lȑ���2:%���-v%��"L]|\{3.�I<q�x��Ģ�_�c��+Wq!jH�$�HC���=�i�/[ڕ���c����d���k��i�b:}l���7i�a��
ܢ.�jq;]M7c:1q�^�ҧ}b�)´�Q�Y�]	�f�l�6X������Ҕ���+ma���o�� L�*��dL�k;")���u�25�=�^N�?aE>���ͺT�����t	��������͡��-]�b㛝s���9��+��
��x���ʌ�\+�8U��Y��t��9}�KW���j{4���=��� �-�����G)��/%B�g�-i]c=_��Jes��p����K%�O2r�Y��T�"t�1��~|�v���'2xEEM9oe�����窰��j�j[m��v�s�r8A�;������&J�:�BT�����ԡH!��A�?h�=a�3�e*h����e��IE����$�_(s)�/����[�USOr\��Y]!HB7z[ת���;��F�j冾�I����l�u3��w.��F��]�nf?Z��> �����`7r�+rƆ�-63x3�'��G�,��c�����k����DI��՟�\#�j�A
Ŕ�� e�([�kV�����#�������dG�tc n����/��ѱV���Y�
����� V�AN�{��n��L�R��F=�{�G'��L�߶@���Z���eZ�-.���C���p���da��S���Z��S�]f��%��&����<�k��{EK}^57^h�ќ�{+r�@�$�BL�a�t��]Ё5pm��°��;׾�aq�es�s�4�2�@���6�T����Ƥ�ꪱ�Fy9�7�?(a���fEȗ���RHߐ���ם��6~#:�5��#Q���)��]5��P���Ͻ�������'��ޜrXMVO�#o����c�¯�BR0�Y�������4��` m�@,��-G�<��t��'�;�����#9��H�U<�Cˌl;���:���T�H<��r�	�Hlڮ(�*at�����7��5��O<�Ub%�&�Q��`S[�E�n�V:��G[�Bh/��grV�������˥�?}����׽S�'f0��Nr����K_;��D�-�48�Q�&G��`$[3n���f�u���I���a枈�K�n�T��2e�"��|���nVP<,��Ŝ�Y�=$��������j~"��Q�.x71>P�2�%E� �Ͼ�e��E�N�x=�Az�{�f��6����-�-�r�����m��y���]	��b$�lZT����T�|��z�,/����#Vź߻.ԙ��`e\�ѷcj7�=%s4U�'��Ҡ:$u�Òw)g:���������]�ᘛH��>��e9@��0ܡA�,ކHv���9p<�~�`��Z0q�l'z���vӕY�$�ejy��Gc������\�ƣ��r76*o��G`�R|�o��<B�����Xk@T�ѮԾ�<7����� M[���J|��v�=�ӏ�M��8�Ή�q0�i���!��g��˸K�&�d�������%�XxpP�)p*���n�3Qt�1��O4+�%��Z��-q�,x����H�P�#Q>��U�9A����
�.k'��h@�'C��k���b/�Y`���RԔ��K�27����K��	�-	���wf��B��j�i0u����E���5`�F���K���RK�3ss��l��7Za�T,�g�wvN�_��n!�B�4L(��.W�/wdz{I1ZN���D�C��*� ��g��� qD��(��<�}ڵ���~.g=�:�������j3�s�'��x��0QnE#���1ސqC���^�.�tiA����&�~���?qY��i�����`�;����ݫ���sw�U5veA�t:���[v3xn���0�;������x�e�پ5�ֲyL�U���]��ۖ_��k�6A<���]��N�/y��{��ɭ� �X��gY���/�+%LSL�.�
�i��0�y��.Q�
}�{+v=̶���ޛ�3�e&��1Ā�;�J���ήs����"�y,+4��f`��g������m6�b��
q�����J�4-��w��&"��.k���
C+s�&>`8�:���%�2H�.ɠ��Fɰ=9���W���#�y�gv���L�j����Z�kk��W|Հ9K~����4����V4�lv�d?Vb��l]��v`w]��Woe�u�7i��^��}f\
��"�ID*m�v��⠵�!WF-�dz/ `�@���;�a�gw�:��T�\ �j���3�e(:����z��ѿ�/�eu"InIhj�b>�2���x������qG~ya�2��4�bcf������%l�^����9	�à}n��Qo��B8�|,����~;N0��v�R:Cun����/\>��#�*X�Lq���:�8�w᫃�b��JN[�>Q������+�E𗝰�Bg�����4E�s�|�8�L��TÒ���B�[i�#��]�kP�n��I�(�-�{+aE�0=n�T���kr⡒���v!,�c49��ށ	���\a�С!1��}�CW-n�ݼ3���p=3�ڕ���q��.���%�6s+�����Np>����":	c$L�U�'���ȹg]b��}�{��Q2����#�3�#`�RTt:S"㓕oX=gK^�~�V�T�r�JD,�i";1�^,ߒY��#�@�~̓����nCIhh�)'`�Zc�����7Z ZA��$z;�H�D���>�=�S]���ܤmR�s������8f�н��s���I
Hy5&�&�;W�-FٸӓlX�@6#���K?�0y��g��u�1��?�V��[jUVe'm�q+� ��P�Ҥ�
?e�P���\7�5":�O}�Չ���;���|��@zU)^8g�H�2��ʞ���6���̧Pf���a��\�NZ# P��tiO&��c���GLC6XV�[��'��L���H<�n���"�8�Z�d
� �{ J��@HCS,?�:*}�%w9/��G�Sn��z�[��L(ƅ.5� ���T_p����z!�����x~D>��{����.��W�����[v��7��v�đn~O���8�1�;Z�q�_2C�����\��1\đ���ڒ=ȧ�n���χ�:nފ$̱��ٙUO�2����"ϲ�����u�
�#����d��!l��
ǐ�Y��jd�,����~�n>�L6%m;CJB�E�Tw�,�&J�W���ʫ-��ץv����B_z���5|�����6�ըX����(���t�A�U�&�_�c�ل��������_��5�ep��Ŷ�� �o_�0՛}���&n�|sw�Y�E�u_�ϼa"g�U����w���.On���j�E���00e#[�~{�5�@�G��m�FUT
S��Ç�p_���4)�����še��uuf�T�/���D ��8����Y3�p:?���o��A���>�)k�A��:��Z�?���0�\�`�lIRs�:��\�S��SQ�3�+�����]�d"s�?�)�ղ�[<)��l�J�����6Y�sX����n�&���=@T��:=;�߻_'k�a��e\��
B��i"�}�e����y�]U���Y�+�rQpF�e�G�)�~C�o_Ⓡ�p������o��X�q(�:8�%�^��Uu��R�`.��s��J8m8�L�UW�7d^U��<e�����N6�Ǟsܢzׄ��g��V������������[ԏ���NTn��nK�Ɋ�pʖcu����e'�>��͢&�㹈^G ��B�d���Z�JÕ?���~���NU�oR��7k���Ro��>bx�k�l�(w���!�H�a꠨�y/�&n��� ��+�ܻ#Ђ~#�OF���`[�ccCW�&K�ݱٙ�[8/�J�e��[tlJ*���~[�qg�9�17�_2)p-�@6��T5/j\��b`p��˹5۬������S�h���.HƲ����R%_IvH�٪6R�n�NK�r:NaKq����P~ʜa�V]S��$��hb[���h��H`?H��b�fގ�'Ϡ�����;y�0�o�l:��:鞊T�^ŵ�)�����|϶ޙS)�`��k�\��S/3ܤ�Jd^�H]Z�Q�I���v^(�K�:�v�aNR�\�s��!}^�𭧾p@�.9T='k(�Q��*�j�z�X�@��E�r�z�9;4��Ҳ�Ր(��Н�d��^W����~'!+��N�)���'#�á�D�Z�p�Q�^.�]xz�q$5J���ڇ�1��4(Ѯc'�6�>�{,�ZJ�o�$R5�Э)��1��������#m�Sa/}�r�UJ��1�[$��Ǽ�S̼�V�����T�L��n�N�ā� ����tG�X�й�˧��7*��++g{u�a��8���	#�fG�N\0�ɔ��z`s$����,�U��o"1yR?
��J
�W+�<*�Z20�ک�=?塀���-���e�ڍ���Ȇ��s��^B��jҳ;�r�a�G�}��q�ړm\㺛PU<���~:������&&��0O������i~$`hZ	R
3W9�,z+t.�L��kdz2�~��I���e�WW��!%��8����&��{�o*���^��e	��!0Y�;���/��_}���Bg��BIv[�DM�^�R\�JDMj��wI��y�i������ G�튿E���
��5(��q�{;Yw��6��=R�(7�X�c������:��`h8u9�i.�M�+���3wN ���L��Z�������o��g�d$��]��=������.Y���)�sꁙ�%S�l�����%��v��J�-4���|-V<B<��d�Cڟ�=r1�Њ�w�_���y��?0�9�˳�n���N��U
���^Q�� �G^�%�8]�k��a�ԔC���6>�%��vq|!��"?��2���?���y����_��Lq��^*oP2uN�vuZ󄞹2�i��0ܲ5�l��(�J��C��
�)	��렀�,,�\��K~h�;��,��VT�=J��дM�����Yq����ʙ�.���"�c>�%�5&?����N/I���-�r40����Q�$b#�6��%CDyDlf�L�9�t���sh~��ث{����I�?-5�Eu�
�Q8�y� !�� jM�~��J�R��7���*������ 3:�v���F��ӈA˰1!:�{;��z:�˟����6�<=n3���P��f�$�'b�f>"0�nF �[� 0�~���coM��B3�~`�_x�o�Kk�5�j
/v3*!��<L�)	�e/B���i>4̂6�쟆�[X�qy��aܾ&*u�N��p�R�!'i2#aƛ{��a�{�"��hV1���S���?b�M�	��~�m71A���:���)�߅���h���ЩPQ ͨH�	v,��{��5T��}�D��Z[c9�{�u�5]�e!���aXH�>�c�0NᘾkU3V���_�oK���АU����[��c�����7d18�#�-u^��yEU+���1��i
��U�#��b^��G(	d�ص���̱D~��0��N۔4�e��﨣h����!�V��.�y4��N;�%Д��72w���W�۽��=Vscth�6���2IY�]�=����j��r��\�#� �`��	
(��9*��-���зw#=�R��R��'�:����^Ru*�����-;[߈�1-hJ���rj=�#!��ǀiZLgv�좄ܓ@�N.&G� �
|U?�/�R�M��S���cdg���]6�ϩ0i�o4B�t�=��P�,D�j̞`�EX(۳���j4fҼ�F�ΏnK5§�j$+6����e�dV�Mxlw�[�܆{��,�V�m�i �:>��l�&rG����~�uc���"]��/��X�j�fZ����j�������\$I˄���8�F�y����G�Y��f��d���-վ!�g8���'&m�+~xxJ�~���<�T2d=�Flt���3�����Ƴ��%(ٹ��@�]���\�HN�~+�ó�R��2?"�ڌk����aK�w��#6����fXd�og���g7T.!=@���}�]r�(�G��1̹�����K_;*�um_#�sd/0P������Y�&uV�i9��_X}�ui�<]���!bA�� ��Y���.����O����cÑ���f�*]��)� V�B�����[�i& z��q�cu�4]�Q���0Ȱm�o�|U�G[��eh�=�\��S;�OoÔS�B�����Tm��S����^`��[N��$s��r|m�I��#��'!��'e.-#eH���}�d)�6���PR�t�$��r�.��HʸfQ/��C\���Q�	��& V�*��mB���Kbu�r�}}�56�,&9_��e�.�2® �p�0�-ڑ��)h<��Z:Ʉ��1g��͋�$�T�n��!��畤	��?��+��oD�kp\R�nlj�VL��S���I6pGk�����KA��e���A�f��K7gn��%?e6w;������8�U<��!2{�|Y�W�O�0����ڽ)1�?�Fc�|�jPgٗ>���䤦6*���K:�mOϡ����!U�n�3�1�-h�9ؘi���Z�t��<Y���^]W��\���ĕ>&~K��R���*�6VE�i{r��l�)Z~�OL� ($�'�!�7T�ʩ���8�m5��A.��(V���-;��{�K��!�*�KXV�ۂ�5D�f8�d�ώ�i�V��k���pa.}��H����FmsL���g/1���HC�4��N���,]��:� ��s*�,�o�۳^�h�i��U�]XJlc|��?�\��3
H���7�}��,�ݙ�����\'��n�8�ݻ!X!0G����w5,H8zO�b}�xJ�G2t��';�H��Ķ��M�������V���!��#AhfSV��ٷ͢b���`A��	l�
C���-����uۜ��=�L�Ψ��޲\��f�U��̋���ʩ�}�!�F�Fm� �2*���o#�f��;���s}tq�Ee���f�V���M����T�^����}����=��u����1"p��|�ߗ0���',��W]�J[�j%�Y"&~�]���	y��ф�^>x��u��Q,�zf�,hht�,�~�E�8X�u�.�ɢ�[��>�pL����C<`I��fN��ǔ.�P�]�bTja����b#��/;S8����y��a߀�3&�!5g���3:�i�}mvb����ܒ=75�u�	A�jh(:�;3�dhR�:������W��5O�Dύ׸}�{]ۄ�ʯՐb�%�@&k��Ⱦ���Bm�ځ�猠!�B�;Pzz�vࡷ�ӄw��XT�p����.�W�Z,��Y��G�)7K�q�����;W�;���n78��k��;$�$m�ĐiX���ӓ%Ȕ�J�xvsT�B8��vZ��͍�˲�d9�n�"�d�y��p���߼��JAB�)}�� �SAR��߶���#�pn�1�0�P�z����aWT�m���={n,3�ǆʹ{+�}��΁���ʴ�,:I�*�BƯP<��(hc܀������� ��b��ds��5��P�S�x�f�k{�	�K��B|+��̀?ZP�_e7W�#��9�~݇������'���<��ۀ�'���j�w,^������3��^�]���
|t%E���B�]�ُ�P��#�No�IIv�n��P]ڙnX�3��扼ȩV���d�a��9*�h�5U��_(3$�ݑA�J0�[�}�	M��'O+��rp�2M��/l�E�Bp]j�1)ݹ���<e>���8��T䖠�M���G���M)L�m!�!���!s��X���V��MK�Yw`	�1@�7α�{Q	��Ic�A��Hu��ǯ���ӛp�!��8 �`�z=k�8xN�3 x��0�����H��[m�d��0�+�I(G�֋�I�Τ��V�@�ü�ޗ�8��A7X\ͷ
j:�10i����SB�A��h�.6{�N|w�{_d.��Q�b9�+;�?����W'r�����JĞ��`W�3SDMk^@@L�K�1�@�!8R�ޮ��;�n�Rr��C�3t^7�'�v���;2��^Ni����&zw��u����Cq���Q̿�Ͱ����-���H�z�&�{p�x�Z��2ޚ=hx� n��7S[������d\�Ks�|�L���Of�}uG�����%N3��$~�80����&��Ҧ��a!k�+F��'�!�N��:�)g��tQ��
�:���.�e�u�{�����x���	3
_� ]�gQ��w�gՃ J\xC���D��&p�<e��ۻc��)���y���'զ&r��![$��.N��n�j!t!|�/�px��e*�1�����p]�d�d�F����n�S\��������+V��������ռ���˜�����!#�C��+�V5��cBP�Q~�`�]��hf?�_B�8�����E�i�܁(xS'D�.����!~��$8�̟n��w2⸙
��Tz,<wn[)3����h��'��SL��Ӛ0P���|���)���ݷ}�~	�NC�x��g��7n�j��90���*��@
9��ʇ �']�2��J�$-<�m���DW2ZJB���'�����;�_�Ȗ"��t�Y�k�蛂�Xވ��|�ŷl'����Q�
H$�����r��[6m�Mp����=�	��P#�]I�P@�}��j D��Y�i�~��7=�J1aB(t�K3�&6��B�B6ETnU�Qgп�K�#�,e_>���Fc	#��ގ zG�f	���C�recq_�3�����)0zg�6c��%B`��������G�rU̗w���%'~��$w�F*Ԕ;�Fd��U���Ⱙ\o�Ge7;�)��MB��y}}N�=�I頻� �O�<n�̹}f^�Ǌ�j>���a���n�B0aߡ�Ӹ{�c
��J*<���v�m��Jx����E�E�}vl��"4��5$FH���[�SRk���Λ�-�����rx>�"fID�����,Ԝ��  p�;ڟ[�r0Nd��e�jqĀ��x�|�֝�fJ���=Dt��ܐ�F�a��S��z]臄]B�w�����{#��R���鬸?Yy��<[�y��Z>6}�R���"�:�U�ُ�~�	���Ը�5�/���0���3�I��hb7#45{!+̷sU&��Fb�s#�]'?]�=fJ��>Z1.������U�'���S�A���ƫ&���ԣ�k�{,� �Nܻ����������V� ��3݋�>��q�D�� r��I6^��	�2K�,�쇙�C�>��37��%ǡx���U��z����%!.��ٰ A?znM�ȧ�E��P���@�c�����_5d��Գ��e�"�z�ݳ�ʼ:.��ɰ��f�2TXa�P��yb`�P)_��h�@�҄�1� iO���cf�R�e���CD�*�Уݚ� ��s���b��R(c-a�w��Ş9�9��'��ˊ1�LM.`��?��<����0��\��PT����V=�0�.��f	#�|ޗ�t��@�?.i��1�WP����$Zbt0���O��&���Q(@�XyU�H�����m�)��C���o)�x���,�P5�ɉ���T�E|�>����V@Kr�9&yB�,����/�P�k���.�]F�#m��;,�����imIW-���t;��2ټo�]�xG�XѸ��2�;%������4*3����p�s�t�q��K�I��������c��w[�~&g���d>YX�,)%�(oX^/eE;"�*�m���<9%��F�j&O��Hdy��W��1Y�l4��8��x<����`î����_��L���%��V�2�w5��{��nF����G��C�;�� �kxfEA6����?�1�LbC�y��[���w��'D8%��`~����Ȱ����J��*&^3r��-ߘШ.����C�vc����ç��i���t<���l� C�g�+��\�foVA�Ón���[��{[����Y�o����L��+�M�X]��(V����k]�g �l=$�����_���d��I�2��П�� ��s�D۾��̲\O{��i���� Nq��I����|�3����䚵�����+�z+�[���\]c����u�K�*���4ܜ}�G"r&ӆ�B�CQA��&��:g�38���9Ж�h�"��y���Z����L��Uw����b��D�r�=y�ɺ�b��Z$\��+WްՁC��0屈��<!CAȔ`�3 ��,�o�"^,6�S��2
��l�hң�������!�@�䓨�obhIo��|cς�(\������nC�8g�t>�Cn�XZ䖁z"���jyWv� Ǥ��cj���VY����Db5��T� h�ΫL���	}�qrc#���8#��$�q�i��wc�O#1�$&.F�l�hAu��/��I�3@]�D-3�ߔ�t=3&�=.���#U�\�q���� bd�f� ڔ��ɱ�g(��t���E뽭�a�vzK,N�;=��g�у�s��W���0����~��f2�|����HS� �3�� 5Α$p&���l�et�� tc"�疦ڧ��%_m�d6��i�>�[U��n"�2�(�ʅ�Ɯ����E�y���˓��^3t��]�~��'�Ы"��ͥJ"�\�������~��]����n�W��L1�s��5�xM�Il��І�7���`j�+o�Zx;|��L�����)"�ng�}ҹ��H�t]/M��I;;���@�������?���R�E_�-@ 5���.��?�ױ
�$�6$#k�D^B9�M��˯����"4��H�
9w?5�����X�n��Y�W��C��K.�II��ǭ��ݵ 8��yl<?�'���:0NW`X+�,�ؿD�]�g��!9� +t,�A~��R�\���2c�g�J�ܱr�|y"6�0�^#~q�H�_������ӄ�-XsAC5K�1tH3ݻ����)�g%�pm�i�H���@^��x���+c%Τ8�u�����Z�[<����5G&觃c_�jLD�ؚ�|<�Qߚ���`$<���]r�]O�[C�ٶH ��Z�+(+���FJ���`�h���s����D�K�� �FKD��lAn�
�/%�Ȥ7�A�i.8��Bq�!��͡�N�"���Z�_}1]4GȞ
4Ռ�W�[F��Ҡ|�GH��e���r��cˣJ�D*��h�����X�<I��T��0'؈9ڊ����;J��� :�~���Hh���3�"�^V���s!_3Ha<�9�b
0*e�OP��+u�	�^@ -�	w,;Q��.�OeltJ)��-ڙ�h�-g�+���X`�j��㱿0����:3����q�[k"������Ggs����-��y��XԺ�����D��9� �D�w���<5w9�n�Ht��y��1�tC̕�3a�b|�q�ث��HF6ޜy�MҊ#)�Q�XG�����w����U#U6M[��-�s4�3O'.����BX�������%�;�x����0"��U�	h�$%�}ڸ���{�5w6�1���޺%_}%���T��N�2K�K�^Gg29*��=&+��v�{�̼"7~��l��<�+F{!�z��ǯ�痚�(b�ӭ�|�Q���qQ�S�m,Z�ګލq�.w�L�/�1ԯL��~����6pq=!�-5gBA�7�-d+/����^�Ň�,�P�`ӿ��T�/��0}�d�����ÈÖ�������IP���#��H?H�\n[�h��a~�>�d�p/��_?>�֙:�^�г��f}a�nk�[�H��z�Yp@D߇�M�'.�0A����o���%"<r�j[��&P�S雳tH/�������b5r����o&�	v��T�CV	�8:W�p��6�/
$��MB�sdQ���j3�"�J��9���p������8�J}����n�!�8��i�f��rN,��ݸ��V_|�%}��_²�
@'� *l������B*r�����dO���~�Hg��. � ����br�~(3��m���o��]T0t� l=���~���\7K�6�iTA�^�t���9��Ie�H�f�tɛl�1���PT M�U�@qc_��q����2� ��(����v���gz�DU:��P6r�2����O��(L�A�wh��bP	�skx��خ��2h}7$��rb_,��?��������`K!Y�����\�0��_,I���:hW��vR�o�=��ӎG[��j�S�c#B��0)�ڟ���[���!����"�?����x����4\%'h$z���`�C7U��8��a�$�'#�_��P�W�e7|qg���1�#��O�3F)�ښi�T�0��g~���:�c�K_F0�[�o�&�oigӼ����0�o]�?	���`�M� j'�ϭ`1܆2/ڞةW��P���+�������k�īxک`ym�� ��u�W)�W;-"�����w�P%��������|�}��6:=�!"ά3�cI�9�����kkH[ւi'�x�3��W{V��jC�8�L�]t-œ��4l����S�:������e?�|[��K�\[�C?V��:'	Ύ� -��\�"����UG��{��IDr���������~r\�Ђ��W���5l�G�7�����4�̲`OQb�s���i]���m[��J������j4^I�&�hNJ
�F�����]G��A:�T���&%X����~��D� @t^��x�G[��qPDR,�
�Pwr�q�Ao|/�B��/��d/�����"\A<�A3O�'v �]`Ӆ{���gDN6��8K͊�6��s�LA`�$g��
)*��F/�g�S=��X�>o`��T�XB�T���Vs�u�����^&�U��� ��Z%�1E��[�,`���g���٧l���i��xgC�c��s�tĔ��B�D��6�I�3�!�N�ϩ�2V�WA��-�k��-0Dl�ٷ.���)�ގ�#:y�7�Ϟ��ҙ`�m��/�?&�^vz���!/�e�^0�*c��"Lq���/80O~�Z�z�P���Rb7/��n~',�А}�Z63;5�u�&wP�\�ϲ3u�,���_]p�s���{y�J����72�ϲ:�fC 
��F���jQ����K=\/|�Z�%�h�#}���<�	EJ��t�]&����T�Bv�S�Q�G�w��|��Ө�r8K,^��� I�3RS� �I=�}��(����[k�z�)")������	��c[?[�)�T��'�寨A���P��=����έ(I��R�nn��*[$��w^���{
܀�<= �؊�j֑��~rf��3~����b�Pl,��k��}M
=GۘB�וO����մIJʭW�g��b ���w�圞�+�D0��p��(�3�<�t�k�X&�7�ۈn��dwK�����*i8Fw�ɥ�G���a�"}&#Z��Ώ=��?��P4�u/�Q�5���y���ĸ��!�BY��(�2Q�����l���|*J���k�;"����P����(?\��=83-2h$�ύ��|���;�|^��<<���5$�<?2G�R�P؄�<?,������̪;���ת�n�����9�����L�fё9�����~ ���v���ɡ@t���8�<n,]��D�H��ʈ{ʕ��.�O�i]b#z\|�)~�fr�k�h,��g3 �>I��x��G�e�l3j�MVD�,���z� ث)�f�����>	&qh��KnZ��P>�5}��)�3��S"�M�b���Q����H���G?�C���@�أѼ5�b�ī�y�+E�b`��L��z.TN?#���D@ae�6y�d\5�T͐Y��n�jo!�f�R6�}�<Pt�I�Tj	�E� ���FH�|x����q�Ǫ��/�Yԇ��B����9�1a���&I�l���z~���g2��!�.�[_?	ƅ�Le�۸���NX� O�c$m��I
�����"~<Bᤝ�)���d}�t�;���`�.	�fH�92CE�v�k�l�6�$�	x��;E�&P�ճD�Uo쫯���2��91Q�����_8����TI|�aq˻[���]$�R҂�L�zپ�f�ôU(��|�7��tR����UX�������� �
��\�����x�����&{����g-W���8z�]�h��,�VhI��g�����.�kk�?N"�k��I@���ɗ.'W�WG���z��e�Y\�n���3���.%*C�˔r[�0�!y���9���{�df�ۦ�G ���Kyq��,�}�:M���ҵ�{�&=@�G{/T�%٠�"�pc�Vɿ�� �����ѽ�����{=�M[B%/��9)M&4�*��>m`��j�g��N��Z�`���iBT���0p�kaN�'��r��BڝEzӈ�1�A��ݬ�̔�eڄ򊲁��Z@�,�MD5�~i0hsw$� ��^���O.�a��@&�]̔��U����R˫[<��aK�CN^[u2�4 ��5����Ğ�P��uZ5��@R�I�ы��S�7���U�7DK�����UD ��\���t�)|p�4�Vd{�:l;"�����Ǫꢐ�5g��B5w��lA��1N"s��)���������PZ;߯0�0�w�VY�_��؏JQN,0u7�_t�w���|p�P��l]-�qi٫�4��`��%�4�@,b�����|;U�fg�� �U%��v�`��b�6c�\<y�د���/�1$��#L��/n	X��:3[�E��9_�\�I����(��t����0�N�e�7�{���lo����n�NL;�}�arN����$L!�@�9K+�[�d(ĥQf2�8�1�#6���Mg&���Ϻ5�����I�_ѩ�_#T�є�F1๶i��ۂ��j�ԆS��ܭ4�vsUK��C<�r�<G�o��-G������ ��m*E��/a�#�G4톃$o�?L���'�
Ҏ�^�U���� �"���p'��Щ�y�aa�*�Dl��\�8%�����ԇ�s��l$����?�1#�,"�c+�$(����w�Y�tGm�oPaGe�V=���a9��@`�aì���>�x,o~��$�0�^!�F8RI���t���C�}��}m�˒B�s�Җx(���F�Ӌ��.���`t2�3��x̬q�t{��.�j����|��,�;D0O�Ʒ"�a�8��.�ij�>Wzm�9�����a�+���,��`�0ç����!>!�\�E�!�Wd_��e �M�v���L�rD�g�)�H�44Qމ�SG�:�+6J���u�=Zd���~2���_2�8����78H
�HKi���c��=���Vڷ&�R9���Q��ߔ����>^_�? u�K���i@���,z��@4{�]*	W�3�祖���ŏ��:�M��X*[�/��:�ש�}���h�$ٝ���xt��˯eM��Z��&���#n��7��d�ښE*	6P���A�VD�tm�~H���Qɥ8J#�G|�:A��î<�He@�H��	�lӶ�{.m��Σ6+�I[�?��LkzEiˣ��&�݁�BҽV�з���E�;��P���=�GQ�����漆~U�����<rCg�}�_A9��shP�ǳ-�n+��-�P��
�W� ��7%G0;/�G-�p��������V昬�#b�3P3}��8\��y���K�s�u` ���Aft�Kc{*�:���|Y�أ��U��߀���(�V^|�a�pd#���AsMi]���+���d�p/���Q��e�MeӀ�
=�]!� �(��*��J���
����Ϝ	\2<k��; ]gzX�g�ح�O}e쾓o�d�%Q-�ts�]����X�1��@p���[KB���Q��jT��rɎ����tI�,��}���ё=֑I&Ǡw�'	$��hZÚF$/��~r���#�w�v9�LTa�0���\r��ޅ_��8��=���f��p�i5������U����t�U��!M�{�X�C���1�+��j<���x�F������R��	5ң���΀8��@P
lE��9D�w��� ��Uq�5�_tbk�~�O-��R�|cEx��̙'�W�W��uxOT�5`�m��-��T}�hmN����;|�nn�m<c�!v�4�Hu�oR��u�.��1u��&����m!N����d��`��x�>��R/�u���-��O�rQ��2��"0&h�P�:$����Pe�F���oj�!������2���G����C�:`�}&��xGS0)ws
��#��S�ty��&I�%a=�P�Ԯ;�a�����=�$��ՏG�h>��MS��4�	�]������M�%/�t�o��8l�:�8P`�*v�r	v��'�<�"K_�ʴ��F�"�sV��5��rYc�u03�Q��,ɭ�)�V,��:�T7N�U2N�1���$�R��K4�d2���P�)���<���,F#�7d�WP��KœLsχu����X^�' l�g������T�df���5BéjJ��
�6�V@G顦�.�T�Ц��_��%�O=P�E�WL�T�ub���+�M���(�s��?M~m;5��{L���<����t�C�CUY�z�8M�r��K&�R��'�T��נ�ڟ�v�V����
����߯<�!_B�K"�����͸�xL߄���Re��b�s����
��A��V�㓺"c1�*�7L����Wԙ��:�%���!ĩ0����)mu�A7J�ۧ��70�7Q%�O1�^:zAE����!��A�t �B^�˗`)�+�?�v�@���K1Fƅ��{+��"\�m$и̧��/�АNB�X9E~�R'Y�"�K�k0-@������E��?��R�N�+ꂭ�����2䩘�q{kM�ը�θ!9ñ}g���j���
7��閱�7 �6˝��	��~ؿ\��x�N�cxL/�
��R�1Б�\�Ҋ��s81�\�����E��a;�����y|g����V/`�1�t��'����skuU�#���o�`m�VPE�@�a�Cjr��rA���n����`��/7�IC�Ɋp`��.\s�3Ð���>9T8[q"=��N���廒�SY���N��J��F�.�"!�f_��B3�oO:*��P5���0'(��#'^�{\��t��p>ɨ�sdn��3�Z/��I�Dm����+�뽥;�OB�B�K&8��Q�&UH�Ź�����w_�3t�s���mb��x ��8�ZB�i�w�Q^�M%/� ��Pih���D��ߺ�A��}]V�	���`�앆�b�� �ux�����0�0ȏ�ĥ$���Y�Ok|u�����<�-�w�oH*�����h����J��9�V9���,y�Rw�z�¿�G��;��h�a�4c`p�s����n�]�H�L�����=x/�c{ H��s�"�����������#��uJ?���Ck^��"Zy�h�z���C��]�g��<��Қ��w#��66�P�$�^��;a�ô�ž�4Q�]-Ϻ^,i��G��?2�� �t�^�
��'Y'������sUAƺ�f�t����!��K�R\j�=Z0ɺ`yI�����y�cz�C�]g�z��8���%��AWcJ�Ծ'�>�C�T��*b��ش'l�3PF(��ә�0�� ��Fji.^,�h�EK���bіk+EN��|��oN;Rg�&���!'<Ȯ��QN�������.zxZӛ������t�lq���ˍɉ��ny�# �������"�i%v_�F�$��x�|�.� ��#B;t���5{�3J�+P)y�ǘ�Z�v����c̲�\�^>�У�	U�}�l#z6/о����B.[�>>�������="�i����J��,�8Օ[R�Sz&0�7#.d�5�>t©�2yG�s��~-�Ec�XuA8�.&�Z��{�I���j] �H���*)��ަ�Ye�bn����[��DV���(��Q@���K�((?����4�=`��-}Gx��M�șC�r��ݢ/ףY?�#���5�iI3@�Z�1�����Vi&kv��+��� �����*_Z񹡨*�� BA���H�%� �76����@e�X'Nw�]H�\��Za�:h0����U���J�+8����b<��a��X��?��eOu���,P%��l������U|���O�ӗXT�W�`p	W���6i!sv4קk�t(��q�Zi�����֮�QB���Oԯ�Ib_�d��Mx��	���nu6��LBq)e�s��x�L5y���h�X��� �*A;�F�--!7�����4r��)���	�)V��*���9�7$��M'}�"�o5嫱�~�����.����}�`�W)�cTf������{CNpa'�jmX$??A@#m�!�^��N��_0&g�.j�����()a��GX���_����x��B�T%x@�Ss-�2sr����{��2����ש�� ����JG��fq���ݜF7�Lbć�3H����~��ju�=���i��Y�IxA ��g��֒��N�/��giށr�p�{�?P-��I0-Ἱ#)�Jŗ֭��~�q0n73n�O�j�;M֚�����I���M�(�J�?�|�ޒW�M�T�oAn�=-���L�?�Sw��$����.^���'��`��<����-�	�T��Tgʴ
P��`�h�7M)�[8����(� %�S�����'A:��THW���
')���=7�!0f��;/�V94.�����1���(�R{j/�Em
R��!A˝�l��
|�pKcҲ�2���萸̝�m�y��ٮ�-�vI2n
ȏ��i۟�DC��
��g ]�{Y+)��QRBq Byw4°y��]a�V�T����Ml�S��OW#d�E��i�=w8���lw���?d�Ŕ�^�dn| i"%�����By�:1G��ծS1۾BYͽ��B�d92�oM3<`�O^��?�:�/�"��BR�݇�@ڦ��P�z�AB�m�}��緧��;�qMl��k�>F��1i����ֵ�X�;5��H�u �et�k ph��s~�]���H�U'bWv�ظ}�V��gl����=�:,�w���Hff٧-�Y����?��c�CU�/�%�Dai�����5��C0���'I�a������l��p|a���~�Ƚ�Ӗ}���K��@5nG�a��T+[-@.w�#pCK�B�����U��/j�[W�'!�b�h�yVF�Oxfy�dtG�&L�GZu���Cd�FO2�)�5k���Su�4�4٫H^L`�*s�����/>p�n�0i�j����q���	������'�v��	�N4h���r�aoO)��߿hFOM���Y��3�`KHL����T�{ޝ�n8���B,f�H}_�9F�]�(�#	w0Z0��1t����s�>K���^�ґ�����KQ7�V�t�7P��Dn�r���p.��B�{K��E$3���l����:��P�� )W�a ����k�T]���|�0�T�ͺ���걷z
��*�>-�y��z��$�
#.t>��;L�O&�[�����c������>��(ʟB�k��k0HZ��a�29��S܂e������d��煨��%�8�d!�(%uXqD[2�|���6���&L*�>�m6?m^��t��G��¹`ښ����I'}os�2S=��R��jyS��Si%�)�A�%JL�G�w����	�%cK��i>���Px-5Q��	��Ĭ�����82��J��(�"�(�(���'mhk�'K&��V�u�M~ �4;��O��
�aC@d����=#�_��U��W���k7�R�C��}�ډH������G;J���D�Z_�D�o�-ʏ�I_�X����Sۅ8��_�l]l��� FY�X�`|�����t���JŽ��t;�$��M�'A(ξy��f2�rŘ�t�t�Q�%� �yϙ�ä�����n�Q�K'	��ٻ�W���}�9,�1���vֈ_A�w ��p�\A/ҝ��~�![�&��h��2��	0�<h�]�${<��ج�^2������y�e����@�-���j���|����"�����3��/&�vm�\D��n��XW���ث>V�/�"޵���n�[�><��$����Ґ���'�	�%�����6�~yD�p���u��Bv�.%��N����<��ſ�G�	Ҡ��JQry:Y^B=_7�wX�~�H�/�2 4_���{)�
1�g9�☜����ۍ�������)���m� �����y�4��7.�iܩ<��w�v'ƺ�3ˬZ^VBwz����{�s6
� �ш�3�Dwe�=�7��p�S*S��T����w��/�iM�鐫k����)�ޗ-�g��	I��E�������F���?��֥��ɕ�.�˘2��rj��� On��_])�ri�,Џ'8�A�ݹ�*�4��1�LC�ԁ[@j��Q����{�&�)�U+�C:(z��!dv��0��o_�e�������ê��i�jo�{��&'�/�Фd��ZJ���j��Y��pI�}_;�
 ��!S�=�S�]�� �.{y��Q�ݎ7]p��WA��KO���d���@F�}�,�JtKx����q�4���]���N�p��č���&���2�XW�gLn_GvR���������/L9�ng,��H=�Z��YJ	��E�&��8	qԔO���9�$��Q�<���Zd�`ٝ�����ε��k�;<Î��%�r�,k�� �|?>+<��d�\ �Zos�hY���i�m#�����T4gf)��0�<�:5�>�����V{@Dka���ܻ��*�)��f�q���jN�W"����́ �S�xi�_"3ɬiH�	���4��y5�]����k��d
aMK��f��ꋜ²��"� `���Ŭ�,�󚭨d�2�Mץr�C!�F��v�c���L��"lU�*�ת�����^��T��>�_D\�L�u��r������u>�v{hǥ�CE���qn�f�Ac�,I�u���P���n@]����oQ����~m��r�oՔ���>JZ�t##,pzKc�����"�U�9��J�8�ΜG�{z�K����Ҳ�
(+��ܝ��JX��~`�����(''�]~?�c�W���Z�Ը���y��q��h	���ᆓ9#U(]s{�얩��S���a��(���0��=�A���N�2Q�e����B���2G���)�r!�Dv��e3EKwY\.�%��Ak�f�7n�6��Ty+Z$rfR���NL�MR���&��YY5�l���_w�B�u�n�j�U��Pݟ��4[iK�!���%�-|j�A���&���i�e�C��3�R3m�<��p:�u�	i������CLY��؋�������<��,2��@<*�"��t��.�nR�@��+���
f��������T��/��6�ŵ
�6�U�j��Lqm!�p���&;M����d8�9��T� 7�AF;fw��q�q��X8��Yjp$��]��|�J��2���b2?�jKx&B���;�R���9p�F�y�F^j��].�VЀ�����C/�P��Y���N�����A�|$$=��1����W�y"\d�Y���N��O���2�{�pH�_�i3���ƛnF�;�ߊ7��2jL�_�l��e�3!Ȃo�GN/��P�}����p0�JnE�SQ�<�y E�?�2�P,��Ln�gD��/z��"�aD�Gtf*`��\�q�����#�'e1�
�ȟ�w�V�#zj2x[��ϣj�8ix�#K�r��ʂ�?(O�z�YF�V�������K�{,Fhޙ�Q�h��g��}NJ�=�C�ÈM|Y����2�i�xU"���?P3�~�
۸�|�ȋaO��~M�׎۞o�>w/�{�Љu{��i�]!)c[A?�����9���[��)����g=3g�c��3�Һ��2:.����StqH i�,��[n���(��A�s�J���:�$�P|<{I%K]�~��N�D�N"���-�^���dkIOei��2g�|�0�*�v����/#0|��2��3s?���.LF,�+��#MV���J���)�F����"❍ء[y7Cn�Vb�7��>������s
�o`vl��{���d*s]+1�Ym��j+�-��w;w[�X3Q�%���N׍��utK���me��Ɲ>�-������Y��D����|H�ǑZ��������\ �(�,�,���I��&
 �AӺ"
��9d�FE�P�N����ķ�/�����184�\���:y�5P)p]�*2��0�R��i�+�3�6�C�T�V��O�rM�	������.:�Z�.���e�<��p`�3AU!�H<q}��HX/&",��I���=*rޝ��NO�6��"5O�b_�F��
;Y�7RgA�i��ŬDf���`h�y��X��ͤ&��.z0��tN�zo{�>�Z\�T�;&�<���`��֝(-b�,��sU�s ������@���*�֋��E�;X�v	+���R0�sk��b���6� �t���^l��Y��,y������b�%��_4�<�gE�6�+�(;>���I�gohr2�|����M���$:�T� =�-�J)<�4�Z���ǁ�TbT,�����q!>%?+�,V�O��X@��)�0qW͍�~���M��+.�X���͸R�/�T{4��,��m���]��D`M��ӌ�YL�z���}���L���L���4�{G��E�<\4Oi����1TJ,.*V����UFo:?>l�;�.��|�趡 ��rɱ^�:�"���B�?�+�s�y_#\{KR|��VAG�{IY�nL�1@?	H�lf�܀���T�����خZ9���fGO�p-w�([5��@rdC{�>8��9��Z�d��[r2}����#T��bh�=k�n�(}��F�����'��n�6~�R�:�#�G9J�C#�
�Oz���I�/3��*Wzks6��r��[���)�PHj$d �o�&w��pnؙkb��!܆5)HN��¦�~6�IȿǬU�2u�\`Q��M��� ����;�����l5���50�����;]�:k8[rT��v����E��O,����M��ʄ��c˹��%�t�}r�8��.�O�j�ǰ�*�EQQ�?ac��Df
���U� Wӆ������@�F �\Ҷ�'���\�l�;��`4ls�	��'�C��)��i�މ�
�l���3+"�t��-��B�U�*~�y���8�.�����PgK�5]C�λ��q�N���&�
�}'�,��W�qAY��1�&�ξ�ݦ[��-����G�NH��Y�.k��0\��ΡtN�F��p�م{�}�`(�.�E,�j��a�E}�)�i�)���=��V���m{͉%��<��r�0m��6ξǁ���\�x�ӒO���L��1�!5���{�M��r5�P�bh�Օ$��x���N�I#y������e�>�j"4ؽFC�(��_o6�����j��������Y���pZ˧}R�T����#���R���f�Fܩ@ͻ�P�Ŝx)=�K��5t�m)�}���@�zŷ��2�*Yښ�5�1����]��(x'�:���&���>	�p���	-�]���>w�4��Ό�21�[��*����,q5h�Y��(hU��S򭌊�W��νK�ÍCz�[��۱fB���J�qI/\^)n��$�S��!��u�)��=�kç�i��ct)��`N��I����� ����6'���'�_��~��f�{ӊB'Kaw\���5w�{�1�eڑ���%RG��;Y_���i{I�N5����;��N��1�)�8N(&tN7��� ��ߚ�ðg���@��8��Od�bѽc7'� �I{�	�:�/��o�~������ӎ.4�#��Qh�ފ�+�c)��8�� ��\+F}x�������
�v���%�������{9s�FKtV� 7���1I�Rh��8އ�K�V~�6���v.�A@�|/~���X��&Y#�C������I��\t��f��@�b"���j��%D׊��AnS�*^SP�Yw<���?�lA�1�Ϛ_����C�铌�LTk��m���m�9b�4� �"
c6غ�js���q��l��Q�sY�"ẚcGq�P��Zmr�����=���c���ֈ�����}}N�hF}�u�1��o��̊+�;X����O�n�c?��"��$��bE)�G�5�.-��舶�?.�d��.IB�DV��3xq
��}��8��z	YHJYRqѼ� �տm���\ X���8�^�e6 m?$?�IJ���{��h��x\jXń�V]L��'����O�=M���X���e5U�a�&�o�j�Z�J� :Kũ����IK�̔�ZZ��\��O�V�(��9��C��&?-q>�50���+8a��mڃm�B�L\ֈ���aL�ӝ<��|����������_���t��{��*8������t[�$��)�4���A�&�s��c �ZM >x�n�A��S?kߒ#fW?	7���>��&Q�b�\��
��Z�(���
j�C����Wn �`KkP@�5\��*=�M��(I8�����h���Ur����z��P�������΅���ޱoYh�ʊ��]m�Q����d9�q�|z�U:\rF4x���$-���[�jx¤+��cQ?]5hÂ�5i�~:F��U�����ղ�-����Eu�:d��pvA+v�1�C�{���o�6�s�	��sajL��d��gp���_��Vd���Z�1���5?���h���k�ጱ�b.ǧ�f�L��$}|G���z�1߄x�����7��I�&�/p���1�`�xK�<��^���u��ӢY5�_���a6v0'O/"2II�Sa�)�r�W.�͖���d���3!�?��I[���8��t��-��>\����5�W �j�7Qg�
x�6g˦���
�F��Ɋ4<ˡ�<	7V,v�3֊-��q71�9�T��ˊ�m���v�LZ(�{F�(J�$��7�̲��MWdv(��$���9$��z�Y���V��H�����о%X`��_����g"��g֢����x��n�d;My4�-��:\A�'�Q!mI���H���� D3��8l!��b}���M>P��k9�d+�Ĺ�eد{�y���2�F���m��w �D�XF�VC��P�g�5��p�M�����r��ѳ��+��M�^�{��O��'����V�ot��ox����<<��E�V��H�'��8q�ʚ�u���ب�����"�*2\?z�m�V>��"�XU�L�G�Oo��(C����X�'�V�ڤ�w'�f[s��slzu�*N3�↭6����t����W ����ʸ�x\��|��M�l�@�I���ē�G�!��[����>�9�����ui�sZ�2�\��v�RW�������ɹSeMÙ>8��7r��'��l�'�UX7�8�ӕ�������U{y�L�g�E��P}����D�)Xe�3�w~ʝ��	��]��.�Xg�-�M�<l���{�>�37=��Z��N_�?�eS��L�׿d��v�03e�Lr�VM�����xu�X��-�P�{�XK�l:j�F�<�������!:��J���#-no�f=�fK��y��il�z���/��F׏������o�@��<����.��`�^F'��7#ӻ3��@�t[WT5F�Y #����.�$��V0�uX$��Z��-��	,��d&М���b;_�3��Ъd�$��������:	�����V�7%"�r��f��,x&�vK��Ky�i�4+L���U*�yau��%��^�X������:D#�"��L����B@3�&(3��*�~���^�Á�a��G}_OqL��9��pZ�]Q��
*����3WfM�Z�A2,.N ��X��g\�57�H3t��,���P���.v��C�-����A�8�ŷ���y
����݈��tS0��MZ�*s���mߕ�F��]hl���;�ִ@�,�]�b�4�`���S����U�M)�/��J�x�z����8د�Fw0��g�~�^��H}u��8�|��o��6�9+1��_�q5��L��}��3	˿��	n]⿤�up��hmr���j��WX��J�Ń�h�B�B����qr���z���o�JBu\4�/]��k�3�5n.M{螊 ����|�/e1��?^8�����|{�u��n��&�p�գ��V�Y ��.�� q�UX�3�l�c��Q9S�˜���@��>�eh�1E�tE��m�l�1�7�읅S�]�A�"��X�����Jhh2e��<�����$�'�LC;�\���r>�
���|ظ����ɝ���A�DZKl�c����Z��Í+̰�dM�p^IF>�����4^����;Q� ��x�i|�V�Q���k�'���s��Y�p�9�ʰ1��o�Kv�YMQ
?��m�{���{�>�^5��2a���\�(�+�DW�/�X�G[���zrxlr���	�_'���n��I�S��^1�%��z��S�H�B\gQ}���&����/��A7��z�0a��1P�̠��S�D������o��{C��C�#��V)h�Ǧ*��T��'��n�>#����}��oB���FPV�ˆ�.�	���V0M��f�yTP%�[9MTݢ�$)����pj:��i��=��
�C��8�BY=�N�����ME �OZV�&VX����'U�A8�jI�v8�1E�z91�3�7u�x�Σn�-�q�q��?�H���y���>x�jı<�3<��&Y ucL��v��G#�h����a�.2PO˗�0�"q���5e����Ҏ�i��0ւ���S���*���J:�:�ᅢ��h^�"9����ƥg�!8����MfPtl� �,�yD�2�����N���d+2��!�nk��C� �ű\����Y:Z�H� C��X�Q��'|,x~x�����*r`!� ���%wj�"�P���h����v��dz)�S�sF�� ��%��/@��RĔ��Z���c�H��KX��0�p��Y��[�`,� ����?ޥɡ`�t�YAL��l~��4�#m����3z�.���ښ��}��2W″gt�ǲ�� F�a��F3{�!֋��HP���+�V��;㞣��=!����%�K��n^`X��n�j��>š��#`z�E� �X)�#y2^%u�%c$�Dö���)����;�VC�*��l�����<�N�}?gdS��/���m�z[:�rP����5�m�r���.,���D�/��6[��{��&�%�H�����l��h�� 0.����K����������I%-�k�߬��}vbar2���8?�O��VYKV�>.��zk��I>OdEV��G��9��V�����fr�y�8Jg�f?^��#1A��/��g�ǜ�<a��<�~
,��a��Ղ��n�د�Nn�+�1���#��bx���:D��)7ȗ`	bS�˗��b��0Lnm��]H�H`�����S�P����fm�u[�?F���<Ո�u��l�n����u�GSP*�GG~ѭ�� 4v�!��l��4*߶������g�ݓ���Ȫ�xA�l4$#l��k����P��ʋ���9����SbnN���T�mG;���e�nTL�fqH�umy�F�ݣ��H�p��p�n�?�Mm��F�8�e��MJ!�W�cl�SU����U���Ur+P�M\:)�����n��QUcy��M{�I'�r	��is؝�������'erj7Ү�u��������ZߴT%A���WH:R�hs���ss���
��i�hs������U���2�K�2�.]�$��=x.hae�㫪<M�w,���L��:͙=�ƥ��:���o��3v�\��v��2Y�:��S���Φ���b�2��\*s�Owlo�3��U���ڳݒ�,�^�70־1��~Tyzn�S3����E��5�I�Vi��ӡ�X:y��rR��V�gJ���=	X�<<]�0@�­��s��m���j5���cǧ)Of� ��n߃�vd���Z�R�섶�5��I�UZ�NT�\7���w W	R�1�����r�no ��G�"�
��֙~\���S��e�XW�Zp���������;7��1/��1yn�e���@oM	Uԣ���;��s%tM��|��&�/��=�\�԰�%-��	�4>ݳN!(�!w������O��3YtZ��<�m�"�G�R���6�P܁�l�A)W}#����7�Db@�Mh ֕0	1��0\��J!�=F��g�O�3���8-)�4�}�k�1ꊘԉ*�n�N�����#&���F�{G��G���I�xv�ǃ�(�����A�{����(��3�6D ���E��|�!�.( څ��ǩ���ʎ�+��d-&���N�cGȿ��|����4ɠa�\&�bo"��A�SB�N������Z�ޢUE&/���+��1�n%����*�<N���{���i�qT��O���ė^��Aư�>:q�GZI����j?i�ŎF�9�E�ת�?�4�@B�aHF<�#���oyW��U��B<��z3�|bv����͙l=��hu��YXr�ڰ�ħ�a
��9��8)�6��l!��˫���w����('����rĚb�I�"������+�_��7;�:��T�ۇ/��Q+�M��8&2'�$�2�����fБ��7E���.'i��E�I�˝*�,��x�g[���#?=�����{�N!��� ;�h��e�܁m�qk#� �B�O�y�L;�oj7 �c����WM���a�)���m�x1@��º(���2�o*v;�}�g<ϕo�5Q$Dn�BS�6�ٳ&(xѝ�M��D����MS�E��/�2��I����C��N�e�/@���a���9���%fX�s�&s�HĹ��1��`�_gR�3�V�ՍS87c[L��d��k=��خn5d����g�c�DV)B��j��!H�/�ީhY��j��Z��7��G�1�Z��lQ|TMO�0-7��k�q�������Ƈ���w�7j��Z�w⟜^ʧC�$���3bG�lR�?�����O=^�*�Oߋg��6y�b+z����<û.���N9I����p�4;�8~�A� �u�y�z6$56���k�c�9@�	�.�)ȼ̲�ئE3�9%����K����n�Dj�������25�wao�Sَ���� t߻}��6��z�T`S{;߸�U�|̾�.�p�����%d��Q�W��"� O��n��+׉��1싎���o�-O�j42�N�Go�bu���5OcG_��r��fr�ݫ�p?��@��J��������i���7˺C���|O��NM	�(�y�)nM�b�U�dSu���4M{�Q��"�fr �}L}��^_�n�CVX�]h5C�?l=�����������d=�0c�j)k3�M��S�Y�����P&�}.I!͆(��a���݅~ЬA_�)�=)>�`�;
�H�
���.�}B6�Ά�H�0x�6a�7rƴs�9=;E;�K�$2����p���
Is���P��G�.���d2��]�{X �s�ݧ�bP�8�@hX��y��'��!��;k	�^Ħ̷��,%�J�k�z���A����0g�u
|�	5��������%�wK�����^�s�[���cC2�v��날�"��� '�=�1_l�[b���K`�P��I���n?�����P	�t�4/>�F�o_��-0|�%4�}��I
t";D%�E�t A�q+��Mǈ��P��D�o1U�<5yI+��Q��o3���B�ߔ[�In���{섑$ݮM>��>����.e���a+P���q4�+�D�h��8��4$|\�v�Bhv-}h�<Jfr�j��~3E�.'�kș�sM��1�/�%ɷ��\J�6q-�t�W쳭ۃOǗ�q
. ���aE����Vo��O���I$*)�wb���\��$��nQ�-z�} F�V�fKB�h��vp�1nh�x�q�1[����� ���q	#��te>%Mpʔ`K��c��J��>����6�[O1Ei��:��9)�N�爡�~�Z������ �Uc_=�X�pd
�<fP�4��~�ϫ��7��ɰ�
���b�²�ǐd�i<}�q'�`��!_H%\*�07F�� ��6���Л��{��5֍�����Z��4�TM��f!�I��Z�jأ"�֌��+3_���Ђ#�q�4hdQ�Q�VS�&&*Y�QL�>A��c���6 ����aH��J���<�-�9��F�aJ�=�fו,��H�1�{p���b�$
e�K�Tu�p~R�QE�VY��P�+�\���.����k�w4��u�c��^W.U�$2��[��Yb����g���Kk.V�2p\���tJۍ��g{0��\��'<7� ���LN׍��£��w!�H6nQ��:}�[�/�8sN]R�f���5�b[��j��f�(����	^��0�?�~U�\��c����Wr���4	9����ӿ��X͟���o��=w�����@�3�~[tz��C�69�E���tP-.8�M['�d�Mcx����ϗeq�i�-)F������C�F?���D'*�_J�(�dc�*� �a���{��tq7\P}�����!�e|�&oɼ���{�"�����?�/蠍�ŏv�/�1�4�Sկ#P���������m�T��}S�Z&3;��q�}y�!i��k6�Q���z����>�E�3F��z%l&3���(p��G�&��̀iWhU�	��d�����d�tlDyKyAo�y��]��4��Og�<�U:v(9�Q�).��k���s�'�'��`;b(w}�Y�#_��g��̦]2*��V{�l<��:�6�%�����|ΟZx`�	=s���uK�׿�#�C��S>w}��p��V�U �r������֙�0��$���n�EL������x�[z{��=���.�p,X����	n��8n?aߏg<�u�.�5ۀ��p�3�vM\�@��J'���S��ʨ�-�E�Ý��H�M��PT��	�C9���:ə��v�h�;B0�H����c�� ��3΁��^����՛M�{�#���@k��������M�?�`'��w���$ma�cƢ%U&�YD����������.�sz+'Ja�5f��!��+���h)K����2����h ��s��#a��
e�5mU�Ǧ����M��&�\�\�#�Q�b����Qg]|ͣR��uHV�2f��4J�V빖"��_�2���@�6_H��7g]��J�3���2�^神�t+Y��7"�4�H�pE�����I�6�����.'詥�z�^���5�;�T�h�~�j���	�d��&+����u���lq� 1��
�'�H=��+�vA��7��W���f/`��X�r�����-Zp|�j��C����:Id4������
��Lx���ɜ��(\�%4Y�nŏ��"mJ&;Mg�{���T��)�ISCuf>�K��y�Sᵷ7
j�|:��ܺ���N;f�` �5q�	��̯u#�9� �!X�����W%g�9^�\�&����Z'
��#n����hS�@q�D�1�r��J{=��`�(ػ]�����?�;�|�J�ܰ����ިC�}�h����w�Q��n���Vk�:Ni��g}����ʸk��|����xq䔲sS ����a���a�����@��'�����������k�=�Y#˛U���C�����_t�%N�!�s�j�瞄���Ҩ*5��N�a�F��n-O����{ʍT��łߦ�������[���чJ��#mR���U��w§O��&p2�ID�d:,��ܫc�}�)RH;�և�pp⊿�R�bۤ0|8f��_-GL������=
����z7@�i��*�Z���$��	����wo�\��z #�r���gMWϭ�F�x�?+S�b�������J��^o���f�O3i��4h�M��\b	�㟡�)�>	޾�q��ݟ��~~L&jXvp��Ct���å
��o-�j��&��U@�c"7e�8�s�`���waI��Z��>��#·�As��B.ӉV����'?D�wL`��@�+���pSw�U���Ӡ,����t����7�}v��r�Ua0n��)30��}�O�5_��N��ݑ�UIq�.�MsT�>��Z(E�-���6�6��H�:P(���T��r��(�I`�z��ռ�Y��$0&ڟ߂��g�Kܚ�lw���"��ɛ��s^��|����cR�b���:��a=�r9^i�
�vl����G��d������/��c8����&�H1jTU �Lȡ��a'r\�r�HhL~_�|�!A�wl4�HW3+����9�b�3�����r�޻��,�����*�<���S �?�~�@����\N�l�_:�^�a�Yڤ4'�0c�y��W���?��.�BCq���*y'	��y2��
��� ��X�M��-^wɖ��𑚱�������ҞsU�
R�`� r}م��g=���k�p��';LA�o��Nٶ�I/����
�+M����Ӄ��5���|)}3���);]�4rh%@9�s��#�ն�n��o�����^9���e�h�g7���w>���i��!�7R�I�!M\O�� �K���C��l&ɱ+�0I��
%���$3p��pA�Rɋ3�F�������:t�c�l nt���e$
�/��N�<�k�G,�OY�.�\	���`�[ϸ��0'3�CD/0}�+e
�꽭P��ѯ�6��<����+qK6��Z��!V5��KΚ���<j))�#�i�ܮ�m*���%bFy!�a�|�1�=jI�����3)�����P��	-�j+�ם��j_�k�&$��Fܝ{�)�63��BZv��C>�g�fJW���eQ���-E�V�t��LqW�Z�v��M�U�C�:���:�!w��Q�Ԏ=�o�:L���.U<bO���`������~�|at�.I��p����~��x]�r>�HcW�i,k�<k�X���McS�C������1����K���ÊO8p&��ՎEE��R�}�q-!���xdF�u��_#H����[R�22<k�m���f���Ԍ�W����nǎ��|"��8|�{��W�x���,�W��]�J��LtNE,O���(���/�|vXǷc\����4�~C�űs���r���t��^d@��5�4���: 4j|�vѭڑ�|�����d��dڴIq+�~�=t�@�,Q߾wc�����Bz�ķ[\͕�!��� ^�r�젔��g����	�$�W`�C������L��<�%oQ7�� �^�K��R������}�������>�ѿ(Ҍ-%n�G��giv?�m.J��X�2ׄ-�sv����ƣ�>+�e�#O����e�v���2�u�qUEj8S�tN���� �
*8��`.�UyG��Ru�=��S>���1Ə�u�X�p�x[������D�X���j�t�g���?�9��v�n�����;��NO��4�K�GaaiF������Gs�<�?�Jd�g���M�f"���v{��9��?�q�iV@^)��Έ.�w+��hVI�υ������7�̽/�����˺{�� d1t����QZ����R
�oY�y�-z���;JD~`�"��m1�3L%��GIV	`�>�2φ[ ��_SQ���H괼��jQ��T��R(Ü��������*�F�	�l���/����'Ɛ�"�\o���P0�=
�]ğK=<H��ʰ�����(P݄(n�����5HG���2*��\W�[�CW�a��=ƽWe�p��Ğ�z��<�[�.�ǞS�-^�b�l�7�pֻ�f�q�i���m(a��H3�0�z��>R\�յ
����#¿��O�C9��ŉ5WBﾣ}'��eB����;�1�=�����C=�j�7ɋ�]��M�<�[���s�_/�����v@�:�y.Jp�rb����M��"}�#�"��ԉ��Ww:7���Q���;Vi8�Q�R�L�Z�Q�$�f��$D�),bmE�0��0p�����R��-ظ��^0���8X+��֤����_D���>�O��Kq�j�5��5��ax;����7��Е���4�Yh�5Y=�ي:Q�"Rt;y�bOK9�$��N������L�����P�4	��,��6q�G����co�� ���2�8b�P�M\���\c.�z�����b���=��r]�5$�p���4�a�N�)`�+�[�x��m��e�r$'�c�J�l�F�;�x��*�(�oPqK��Ғ{ɤ��mA�ָtߣ#���߾�E��]�kg1d�sf�؋�X��xF�D�/��`$t��UJdl�Gʨ���Û��+�V� �)��������/��0��%S��Ԙ�Fo}�j&��KK`g؝i/�����vOR}���ĥr�kf|��p��t���Y�Z�?�幥Ef'��Mv�IG ��c�f�'.����J�NWJ �oO��.��ٵ{��	_R�L�Z�-nd.�*�;�s^J$�\P6�b�9:��������_ oǮ�_o>�*�-s� �z4:
3���.��PW<��M��#� ^�L
V4}X�o)�����Eț�5��.z����<^��8�T ��8�K�/�ؾ��Rx�	3�?:�c������{��C�[�}erᯮ@LlEK9�	�B�E�4û�v>�Z(�,���x��%j?���IZ?�0X^���^"��݃�h)��*Kb	�
7�BI�ǯ���J��륌����|rLq�
��~a�&ٞO`�k˫>+����h���M�Z�O���jc7��ȩ"�z��#�R�Y�x��!�wF}��"��m�\ԍ�:Ƽ���'.���������W���/1�:A'���Q��y�0Shs������\̜��?� ��D�#�6��0�ﻵ�,X����@���v�G�I(J��CX(��#j+����ɔ��N�]��ק(I��"y�>��ɱ�%�*�=�}�տlu�-��Rf��܀�_{��Fhf��͸(�`'zˏ�.�`M�O2$>�ܕW�Ek
�l,��x#<��{���Q>��{�Pl���� ���xi��%-�똰q4�G�G�����v�K��������@ӯ#%U}�.��a�+Df+b_���x5�g���ʸ'�ەת�5�� ��&��'Ro K��M���>���xvJD�l���Pc����e��(-�� ��1�%S���je��[Kc�%%Gg]1-_�ЅM�x~���Dla&�MOuZ#i�=2����%	w��}r����#3�{�^ZNo�y���4U�9����,8oO7����#⢡�$�g��q�lЌ�5��� rM|;�ω<��q�v����^�i��E��*���}6\�F%�јɯ����(�݃CE��Ii� ���FH��3��7�z�3�w��f0N@yS���b!��l�	J��Ӵ#r����Z�;���U>�Z�h���`�b�y�*�\�ԇ#̐���;�l~��/�-��9ڪ
e�zʦ�#���OA��`do�2�y�L_EMZ�y�ȟ..�]B��zJY
�@gN���YL����V'&�t��Qå$X�Y7둡��Q�0MA��JS<����?�qM�ざA�A8�>la2�����"�ɉ��d��d'Gr�}�tQ`�E��t�=�mѧA9[$� ��6�"�qqƒ�L�/�W�����y1P��'w<r�LE����b���"kE���8[�d�D�q>k%i�G���`�]�U䑏�w���ܔo��nA��BK�l�\|a	�5�]�aY���?Q��)�چj'{8���i���f8�ϱ���.���Idd�M��\�{6�y@Pd�T�*�������>��Ɯ�L��Uڻy ��:��<����W�7���5�յ�d�����/V)F�|㮚���Z�j�ECl��ɽuw�,'qA<y��L�.�|�ל�f 1���S�$%/�SxSH���l��@?�Q9�,�4rS�W�b�"8�(�[A�v��P(�3�Ԕ}7sC�'n���e����zsj�|U:~if�,j�.+�SM (S�ݒE�@*�&�n|'G^}�ڥ�D����
f��-D�ԗ6��~5ݐ�#?Co��6ww�e���Fj�_�k�c�00���&ײ�AM�;
ޣ����-�	w4/}�n�����������J�I~/
�/�|G4�����x�&nx�o<'D,�݆�r���Ux:O�����n��Vͼg�K�m��1�O����E%�6jX��
â���O�M �
_�H5��4�_�����Ϸ��OB�>���DT�,�_MF1����2��Z��\�z����Q�ZI2��3�V
 �`�eC��u˖B�cM��|guh
�lҒ��\�Ws�ľޱ��99"�]v��0�ǐ���	��5 �i����{۾k�4|��s�w��
c��v���k{v�8���J�Z�t"h�0t?៑*c��Mu(���������Y��q��.`4��j�-i�q/��re�
��Q�&�g��T�q	ʂ�ȐR���EW��G�&!j� �>���@���m�K��A� i��Vٸ��aBDx�{@�àG��R�P��]�>h4s�����	ajs
>�O�3G�E"�S� 2D����{����ߴf�������m��"��t���s�KW4vL���LS��A�!��.b٭)�ڤݲ%Q�.1|�I����N7ʥ?�#i��AǸI�%�[�:��`��%�����]|�D>y�n�+[��?/����mpaJ��|+���l�c��o'z��궵�<��'�"�:��}�@�ŘZ��L�+(���E�t����C�.��)���������v,�;���0ҡW#͡����s�QХj�9*iF�T�PG[�uy�6�i���w:ZOLG���S��))��c���P*�ծ��/�&L|��K�d˻��v���T�wC?6�r���c����� �P}�
���R?��C�˪�ڼg�	�y�}"<,E��d�|H~����f�=���bLq�Y����4�X:�<U����{�Y�jF�%�?�/!�5��$�������d��:�����Ҳ��V�lf�V��>�+����4�E֪T��,��u��������-�� &$�b(���*R h��p!����+�y�w�*CqA��iAЉ��Y�j��=<����>F�ŘyYh�*됻	�0$���\8_qu�#�-��S��Z*�S�	d���c3"��E�Ĉ��y�C�UI�L%G1&�u>x�-���(`�����0ܡ(��i��^.��J�J&(�eߪU']yŮ8 ������i�?���@�YA���$�h+�P�g��}ZR�NiĚ3y�v!2��lK�+��.3�@�=zAՓCNp�Л_����K?&��[�G�g��F���Ў��	�/f�޹���r����~ <�ƑRX�i��K#�4��ʚ+��vy�Z�|��0)��gq��C
����a�ޛ���4q�pkEJ��[��$�d��{��+��se�<����d�v��� j��u:����Q���%�$���� }P�3��
+�/��-3=8ZI1��j+j���h���[�t�]D�4�����&���ض�K�,0��Cń$0U���nlD���)t'��D�<������f�@���������l�i��O)�{+�dG��C���=t}i?Em?(�k�ה�v4[*Ra��W������{$00�s�[�D�5P<�Ux�C�
�ɹ���1�ƮR��i�t�?������f^���<���a�T#��bQGO�"R�*h��u}�X#����Vi6~o��1�&�[�D���s�� ��-b]���Т�3�F�5y�Q�����}�4U)�A�rat�_��>�/g�4�t\b����2��Ѓ�^��J�~��*.�C�,#[�Ǆϡ5�&"h��\ą��,��������]I<T]�wv���ԇ�C�:p�2��^.3
8��:&Ewˡ���s�&� ���Ҋ�e��և��@3�7e��v�ь\�ų]Y;z����ŰԆ��%�nǥ0?���`��ɼX��g����l��]r�Յ6���ib�2\R������52#�~���UQ����)�)+Q��C\=�)f�)da���.��z��]� �^Z3,�ֺ-�Cݽ�(�	�I -���_t$��{e܀w|��d��>�V�SZ�R�fۑ?V}�ݒʌ� �~�u#��ld�X�[�kC�V�yhZ�����qd�H��G�����չ�����n��~~L�hn�i]�c���0C�g�%���5�iKO�4��k+L;��z���<�I����(�\H��:1en;��n��`�f0��_��<a����N���?���j�K �p���F��ua���U�w?K�RA�������x�.�[�ޗ��%��lD��7\87��XYB
���	0��KL��h��)r����pr ��P�o��
�'�����A���7z��T�I��=8B���� AO������{��B�<s�W��z�A�ҰKhc���K�\`'i8Pz���RZ*��^�*G��g��soz��ߪ��W���k��%��.I�;���A�{烤�~e�����/QH͕�����'�=�� dT�ͥ�����|���
�`X�D��oJ,uҜ0|)��.kdp�פ+%>Zi�rx&�T�6���^W{}m�e���w3�	: "
C�}��b��J� ���M�*��V�n�1-#p�g��G��O j49t����y�6��Ղ7����:EҐ!��L�2��8âM8l*?� Z����A��qS '��<�"����˞��n߽�8σ�6�U�Ц�|�tQ5���z�~dB��O%�#�+�q�|��r���C�ϴ�`���2��6��?kL�i��ƗيS��v8�aK]��3�=rZhڟ�
�J9|�t?�l�R��Y(���P�3'?ܵ�B$"�@g#2S�1x6EAS��;��]����.�/��oK�^Y!�w��9��� �4�[$����^�>1'�(�V��ֆ�1u�[��=x�m�%�̊��aڋ
�Lz+���$�[CmS�7�k6���of��sA�ݍ��;��8ι�����0�;��q���ԧPg[�!՟X�4�1��c�rz�V��y��RO�oA{�,у�!W�O�M�*TԕǘF�� �__Y.���l��j[�χZ%%�l���GAM���D���������*hL�@�F��cu%z�o#Go�9��i)0�7l��`��|iS�-]�$eT!��aX�Ξ"�����&q�:��A����&��o�[��f�q�/�<��A2V���Z]Y~���/>V�U]�>�>,��+�����O�K�_Z������.O?���@	��|�.�t�z�@gCWM7� Ϥ>?QQ�,���iV���p�k��+>�90%W)�6��m��@�I�6�០�e����R\�$����|B�qpea�S՚ 厷^��ig���ߪm�N�Q��mD�P:��Z����9i�~,)!�����J�O1��h���v���|_=C�~��gq���uN���#,��X�S±6�A��5�!�}��F�{9DA��sО�zMO�ō�����:c�o���grU?(�����M>��%�yR��ISX�w��ޯ�"�����Y�����+�&N�I��Y"K/z��������>?�_�3,���FACRF�ɷ�H�jڼ����9�"�g4(�A���7SF&�n0�+��&Ĭ�덚
߅qqN56�L�K�4]�����ݚXl-�Y[���������|�F�(�*;�#���k��hN=��J�B�Z�A�K�PjUE���Wg��d���I	ڀ��/D�G�+�%B'K����hO[q�9��)~�3�y�^�0�r��LY��f��7�6��?vp��$��;�ySʹ)��s�)$�9�o�2 J!�'^���W����3 D����D7R�*[[���s:�������C�B�}�e�*��N�wģ�ڵ7i��[8I�$��Ŧf�������2r@��y��)0�z� "�������>��\�W�TC�̀�hd��/SV�,[=㹑�����T�]`��t�m���y��H�~0�Ջ8%�(R��V��E�m��h�D��7]P��ev�v�	�#��l4��om�S*��ј�s/m�Ng�\U�(ծӾ���k�)��<��t)*ug����@^�!9Kć""�w����mmY�ZN����IZW]�ލ���\�N�)�:�7�":	b���.n.�bq�����.� ��7�q�_%`X8�:zm:��I���������L�aB[l�B�8�S�>��`x�ƥp�E�������:4b}N���ha�����'�!�����(=y"V9�����֛�dA��D8�M	ȿF�/2�,:РTLM %�,��C�����%�#��)�wˁ�mKa�P�P6Aj~P�c�5�4������p��qVk$�:I���� 2�׭��
�g��f|'+r�<s��6�۱W�f�dMS|c����mW����v���*���{��hI���\d����qD�r����n��o���"KÛ�e�v���`��j�d���BS~��ʡQi���y�є�Y����� Kl �.�j�JS�L�ɗ2�}3���]q�B�Fȸ#�����=�Ů��ϻ��O����L�R�G�w�,�S�ynE�Gmu�q]��y��\�n�oI
>��oT嬴�~{c�����_��e��$\3�~�f�J���0�*����[��H�5�\m���>�}y��v����8K��@Q�ۤ�Gg���*�f%�VO�����O�2K0�_dο�ոQU������R9�3�_g��z~P�0\�JBgF&����&ai��
mX�=$
��rWpf�����$IG0X�a֥�W
�b����Am*Uv����9��	
�P6���1$�p'��9�LD;;�U?��h�w!��X ������*{$ӱ ��\=St�B7��|�ϋ]�îɃ�tf�L�ņ�~��HC��t��2��pYmf��k2���E�"��{�D��-�O�.C'`��ǽ?_����n>��'�]xA�^���#�9]2�lS�����
�v�|Ј*��8Wd��$�+� (E��� ������͔!'Rf��7�x�vH�51����e�'#�_?!PxQ4�(�4�6.M�Dmq���?i�m #L�\^������;
{�.�2*J��7%w߹�K`��C� ����=4�+C6�O���VMTV��T� M;��|a{>N-��X�k\�}�e]ǌ�h_y�'��*���u�/�:� �l����@�c�����u'U���  ��𨐠U�-iN�<]�K3���}��!�j	���KA�c��G9�{��콮Y��u�ޖx������4�1�/E-�8yf�i�=��D5��>�"��*+�$z$̆�����[�U�O�\������Ƅ�"�:p��"���ڢ.�3�2�BF7�5�.1H�o�7���:��JGca۶R��7)�U�	<���3H'���d\FX��f��f����xX���"�ʱ!��_����c�_w+��F};6��c_�m:t�����;� �9q#���9��i������ ����� C1x���>l`�<0�?3��\|�;�?��p�s��w��f��ͫ���ю�뎾$l�$�U��}|��Iʢ�i�+7�Ɛ��d�P�������"{�R�_Ǒ"*���o������x�jM�b�����\��Y�
��{"�T��
O�l1�mʒ��"���0*`���pI�s����d�����S �k���A�4���J0�8��t���@K�
!�I���K��r=R� �K�ɘ��V?�j ���С�g[?:��^�����c�3��3����vN� �d�3����k�r^r脺��4(S��υ�o?���@�$����Hm���{��oc����'E��2��`qK2��f|r[.��8�	b�_d.}&c�By���^�^S���d5:=$���)���7��:�d�9�����t�k�z;v�qWy��pϟ�0�q�����DF�WN(���_��T�~~So5��sܮj�6�Yl�5C��l�aya�G����B2�f�L��}VU�H��V�#�}�n���A=� �ҙ���:�@�{6&ύI�q}5��d�w��fqX^���s���T��6ߎ�b9���i���'���і���eH�i��ҩ��ġ�|�n��m����.B���'Ǝ��60�dxI8گXA��d'�RS;�F������k��s��LE�K�nyn���a���b�5m:60��~4�bG�>��=�&�:��S��O��ʶ�cƒq&r�.��5u] ,M����yt��A�*���G�F:Ѣ��{�t�_��)=B{@�����k�d�Ny6��f�9�$l�It2�<���o�訙����9E��N^�����Q~9�tj���"1JD0vK�"�@�`����Z^3�]m�S1	�@��2�y�e���JP�`�Pj�f�rRp!�\�c0j|��:l��Ԥ�pw<��C"V�� |B=���^I.����JWzڪ�8�;��Z쭸�zs	xC�7fH_��)��q���'������[��n�!Wl��:_��֐�#d��ɤ��G#%�"{X����3�V9g���/�����Z�#�;!)_A��v�n\���e 4�a?����$Љ���d:	��ѓ��<ۚ�	=Ыk-���� ź>�Em/�{X3�����KF��E�HU�#�cO����"go�^vK`p��3�I�����z(�	���,q���0Y���'�)�bs�s�x ]p37�J��$a�:y����i�$��f�;�R�X���v3'1w����%�މ�{�LE(̭K�~ʹ6�y�%�g����l��N�c%�ƙ	&M��ҋ�ba%��pBY�ae��Q��W���ˠaκ$��3u�Jxw�ލ��5�7�"�Յ5UG��}����x��p���O"��$�����K�Ӱ����Q_%Z�<N�aAU���$P������8
j��צh�Z5h�M���79!���e�݅ �l}Q5L�հ6�^ 6�������s���f��Tg��-?��>eg��]�s��̚�+���F�xj� �{/��O�謯[���lf�T6ݿK�����#h>�pE˝�#Yq����$Ng.�������	Ĉ9�]O�K{mT�'�rڤ0���A�j��\�+Pڠ������zq𠎐$'�J�e���D�x��A?uW���Z������ry�
0&!�&{2r3��|Ϫ&�s��,�c����{�;n��_T6���3 ��LG^�ӳ�	w��i6����uf������z#ᇀ���3QFgU�
Ӊ� Y s����Up�����=p���d��˃߄{�2 �k!r��[<3��%q��ZBZ�d[ ��@PҺB�������K��>@n�T��d�jl��^�����+aL����<U��o<�~��n����w,t9�J�J�}����rs���>y*�|v����}<�)~�l�Y@Q�(X\�ޝ�/&�U���)ce��e�D�O�Vڭ���8�0��3f��zكh�SUuk��;pJ� |֢��p[wG�t�{!�0�!���!�����Oa@��I��p)8�5�A��"m�XW��kr������9����y���Vy��\ܚE%�Y��>)�V��������]��sXN$B.ݒL�!�Fe�?(}j�p������DSWLD,0�i��}�[?ٻ�ތ!ڵ�P�{�r��n��K��MM	�ur`�g-��6�i�C8�W&9;�Ex�k5���i�ʫt`���b"r�D\�y��VI�!��N��e)�yce�#H������f���~����M�"q�+��*�૟���f,pd���h�]D �B
��7[�k�mW"ޗ��l��Q؎�s�˿����َ^~�M
��o�$��L���	�'�����'���J ���d�6<��¿[��0�)$�>ꦈ��\]�X��A��y�"�}�����6�"8��RX��.�\>��U����'8�Ji7���t~�D}h8�
�X�0�0�،8�v.�d��%�!4h��}4H�=y�*f��َ���M�\����/��b|+�����k˕SD9���a������n�&���0�"�,o}(;q�34ɖO��%fp	��惊���OႎVQE��%�o֢��R���L���r��1#���G?n�q�Z�WJC���u=ٞN�K�b�:U'h��SJ�+'l������0jD���������&��q�|���.�#���ʴL��{b���(��r���?�^e�e?������2E�K��56��V�J���;��h�
\�sz/|D[xE{>y������U�>M�{4 |nڢ��A��d��t�Z�CC�o-����lS'�X,�|�;��������
;w��q9䗧��{+r.���R��P_�٭Q�O�U!·�$�&@��:5��_x��,�W��W"ku���"�XɆH�.�	q�Le,�輠x��Y��D��z��H�<We@��k�d=�-�U�8&D����8|Y�Yn��閄-~-���G���I����[�'@I-�X�hү'���`��ZԊ{Xٱ����
A�L�V�(d�;]�o�an� ��r�U�E�� g+J�O㌳�%3�:q۝�:�{�O� C��:
��Ң@��ݴ��|���'U:y�J���1�� �a��*��-H��~��:���^}��	��fhX�qʱ@�PK6oK�}�
0G=� �6$�:9<�2A]]�����	!K?o�᧫�p]W���F���,��ԥ�H����3�`�[G�\|����y^򑘈���H�u�Ys�zu��v�F#��9�dwҜ?j��=��%_���P�ߩ���U"��HՌ�b��L��+�;��Ӎ_B�`�J������Q�M�����]�]��C�+|�c��e>�ޝd��9�n�kc��sD�Xb_�Fƃ����f=���"wcNc�|�c=ĕ^z�3������S4�������E�,�⍱�V5`EG=���j����n�7k���Bm�Z�z���2->�ǫ�aezL�i8A`���g���A�V��~ z1��V�'( 6������c6�O���&6#��� �����T�� ���h!����գ�n>�.nwUr��\*l�yA�J��ئ�	�J>���o4�=�屝�V��\eۘy�Mm#�?e����,s���D��ʜ�e��vGW�������^��wz�����-t0�8X%�DΥZ�9��-
�wRg��ٱ�ؠ�8��G�y3��Ub�q2��'��T�o�% ���PksXI��IG�{J���B���N:'�"Ն�>D���0�ە���G��A8��T�8;�{���
Nf;aB�-��A���7`���t����a�A@tN2bދjWK��$�%�s�B��N&��kzȬ�d��p��_� ��O����nIT��ʾ�(�N�.�RF( J��F�}?8E��4��{��g߂'p.g���kv�����T����^����L���c^�P�^96�p�3��;A٘ә���u�Җ��5���J���Bt�m���kW�q�.�	Ӫ\�&�zŪ��!�%Z�(�7W����6Bm�@$����l���|q,y�hE3k������ ݧ�-__m�Pn;�߇<�{����.Ŧ�Vw��ܐ�W{Q&�ǧ7Q��H��R�a7E�aX�����0��d]䙫.�{dǲ�Q3@��F�s^���a������"�@�D��4݇zʣ{��@kp�{݇=�:CI����cC���n��zʨ�w>�v50TB����3�S��o����9�{�̄z[�RƝ[%n��h��ƥtЎ���#�#�a�x�|<u�sI��x����=��O/�Q�c��5�b�]��W{���+/�(*�D�w��I�䳾;yVd��wp����0�S��6˔���X��Dd�B���0V.�T���BW�9�����m�e��S�T�.hgJ|���� �A-ж�@f�4U]Ğ>r[�5p�k�Kԥ1Ȼ��]#ck�=+
��:#%�W�)��G1QL�P��%%=���i�4�g�n�tmiJ�欔��[|4˵���U�N�x�qh�@q 	��C��X�Ҋ"�r!���jE������MC��$��rk��("��q���Gq���*�u	��O_e�DwF�bۺ�~G'~�����A�r��z$���(�����R�W�$ �Q
�m�j�~r��+�!I��S���X�*�N��l�j>�!1��@AC�W>	�4���̴�-�����!��b���`��{�A���nrW�4;�^�����J��ӥ��8�o˽t�5��c�t�J^Ӕb�������^�Q��(��<{H������� k�x�$�,�#u���e�4����O]�>�LKpx=��Կ�i<�F�����Jw�]��R��"s1���Ӕ󓀲q"4X;�2�qn�9ڂb�)�����6G�5���Q��څ�9@�~��޷"��E^k!7�IL�`\�̪W�)�4�W�}Ku� ��%,p���K���13��`.�(h�8֨6�ʦb<�qe�-�������`ں��iLE��5�/]ѷ�����	���k٨�m����^���l��A���I8˛j�P�	��z΀��ɡ����������#$͹�P{khe�SS1���>yv4������k�'�}�Zڽڑt4s�q�<����OCX��cգ�5�t�r��L>��4��rt�F: �z}d@FK���m�-���`XG�ә���~���O�Y��`ߜL
g5�i�S�4䠲��r�X_���C�'��ߦJ�.�C;U����w��@E���^|��"ǅD^
���O���o�N��Q��;9@ꐂ[�R��߷o36������@��s���<�oH�v�h��R�c�1�5x�!0��sdȘ��R�Kv+fI]���S��ƧU�߯A�?w""U� ə7�Y��BR��[m�I>�m��()�ׄ$�)-�^��kWO�yi1�:}�SIX�#-ʿ��i��)z牿����@�Gz�����EZ�N:4�M���������M�G��}BdڢyX �Dm��kt�����Uҫ]��������B����çu3��%�$����v_}�c=�^����׵���{��C�����&�\�i!�v!#�c��j (�(��e�YM�
a��3��P�P��Q�1O�C5(��w�(�.��#�?�CBm�u�
e��8s+K�z���}�"���ʻd
h�ͼT�>�7�C�$�" �'Z�H��<%xBTE��42�٬i�����@��t?�Oːf����M�56�(� ӧ�*���mx_�đ[��b\����$L�ԕ&z�~(jX��t$�X!
u�>U�)���	5aj!	�V}5k	(S�!&(��(�%�*��J��v"\RX��fO �cT�!�ҚHQ���Mt���n<���oa
�SL���S�t=�)j�����v�?x�O���e��;�\ �S]_<���o�e�Å.J�Z:�窞s؞��Q-�0(��$P�&�x�#:��֣/�a�s`i����7�!���@�|,�J��>5���%tI�A����los��s��Jh٫�{����A�6�ݏ���8h���?���>n�l��0�utч��+t<���q��E��gQ�+(x�[����?�=�Y��,���<��T�N�6v�e��o��wY2�l�m�3i�W Fr�[̷띲��Px�F�����Aj��t�' �&*�k<?���ã��1@��!k���� ̗�;Ze�%�Қ7�p �+pb'ʙ���. �^�W�`��r��Ē���ő@�"�G	��B��9�x������}�X�VY�����Rr���E81(u�\drD<(q�=Q���2�=�B��#j�-���" 0��0�O��Y��X4x�Mţ�J^�,u)�ME�_��lr�EꢆfH&��.SE��Ea��f��H�������u��h�n�M�nO�	���ӝ�PI�0�&k�ʚ�8(�+�_-I���٩˜�7�]5����V��
��Ȳ�z��|��,�n_� �{�<$s�c�f��ᔖcz"�"�-=������Y�@�r O�� .�׃�ja��8�Q�\�j��	?��	��b��~ߔ�a��3K��벓����W��s��	�sĐ������)�\���O��W����1�w	�H� t5
��!���},���y�a����r���#;T8uhBdq�%(Pp`O9�'j6%�|Q�)��9m��JY�5�>n�LQ�y��v���`K�Lz�؛�\��U	��@*'��
>L�77	9�+��H��t�] 5�Be�@��𚈲�#WF�ϱ��	�~�N�r�����gMˌ��O12k؉�Ԭ��1�Ii���R��د��]�rƾ�n���E�{���	�ll����4�`���S=/�g�|�#8�R1�Ζ�t�Pۥ.��c�x�냫."&Œgk��EAt2�֨��-��OO9Hӷ��v'��{�W(
����D��@��r�X፹���4i��u`��L��p���t��v���)\��3���C�*k�f�T�p���@X��T�5�Tʱ�?��%��9��h��T.�(�I����Ё'ݫ����0���D�`i(�²���N���]��'�+����Ja]we��'���a�j Q��6[��%%�1ޠs7�ty��1�I����!�F�t(�B�752'�9؉m!�A�P��F|b/�Xu�ᩒ���Z:NL�� ��bK�Ma��8N�����^�wp�ww�*t������k	M��KS�f= s��O��4ͷ�C+X��\<��E}/E�'���ڔY4����Tvc�ގrA�ҿ���� \�l�I7�݃��c��\)��0]�iG�����J�S]u�F-pAR�d�Rvg�d@�e��"�o7����Si�k���vV�Ї��r��oچ�����Ω�(�Se��p�
o����{X���;ۛ"����Er�<q���@��q�%��C)��������{�����M�;��O|����4��(x�^�ȥ���]�JΕd��pӪ�L\(��N ��C�Fa��عnd��]gw���t�lЕL ��X<H�vq\J ����4\T�%Ʉi">�=Z�����Y�2�a��:��������﬇	��3=^h�MǛ�b�}L��K˼T��I�]Tc�e�8���D��x��R���������D���1&a�Ü\��T�(������D��{H��w��d/#��]TZ|���ƒ=~����a��i�[��3&�,��m�ɏ^����š��9���#=��Ww�V"I�T˲�fWPXD�!t��ܻ�-�u~�n8h�AN��T�����O����X������(�/� p��^ ��)��*�����@������Ӽ�(���n�+�,���&�p<�س��"%��N���2'0%��7I;�~��}�}6�Û�-���̜Q�� u�:�G�ow�έ�yş~gP� ��Z���G*=t/���W�|ܖU�q�Mψj=ǆSc�t�W��S�')�,��k�X	t�`.��޻m>���i*���ֻ��9U��
�q7R�*��۰��Q>}* "񳞗f�`�]+r���b�O��Z��k��Lۡ������)Ƨӧ��Z�{T2����ҩʜ�OY	c07v���W����>m�r�o@�8&a�Ɉ:-K����s�W�F�E�w*r���9;[Px/N��xv_�!'�� ��}�8�r��A�r���m�!	�^6�v��*�T��6���JV6��.���+{�t2����,Æ�n��T 6������#�1���G���!�f7��\�i:�|�f)�ly�!b�@"���)����e@�/��S����X�Y��)���iI��V�xWQ�9}4` �F� ��0��P�d`&f�+��/V��H���pt�nl����͖i�r��-�;���{WT�%)� $u����U"�qD�l��_�k�L�ِw���i��㪊,9�\�c��YC�y��oK�$&�FsQ�{'"��{��r�E���Ğ3|��W��jy����}�E�%,��ԅ&4?ҹ�2��6�>���D����D[���r!��SyS�G��«|$������#���6`m���bB���C!���聣yE�| 0J�
Hd���h���&K���<������:$u�?�˘�d��@B�kSN���d���/���E���� �0:RpB��rhǁ�[�T�F�A]�H(�d���V H`�_(��8��ý�.���+/�I�SQ�R�)�ݗ��R�!�<�,�j� ������5������@�0�C{\�HD�:2�l���']�gm��W�V��	m~��ϴ��uH��!�5�� jJ�E[�Z����V3�7�Hfj�t�>eRu��x��3�ч�:t���c�2e�F�����#&T���f9��p�N�9�&���(Z�*S�P��d��I�"[�z�Y�^�wuhc(��͋�cT6t@l[��}g�F6\?#���m�@�}�S��~���+����й�Z�s��ާ&���s�tm�2����z)O�S�4)����WF_f��*[���O�#��w��8+j�+�8�'��GG�(�R��.|����Ɖ���`T0�.A�U�Y�%R4=�h��[m:���͹<ש��FQ?�6���)y��̀
ƃ ��V��Α�j?�q9����>��@��sǅ����1�{�����8���96Qd$�P���6F z�`\������U6��W�n�Z�9rn�!�)�.	���q�t����/�N��TQ\|Z~>�2|!��|t]h��=�;��Цǒ�J����=!h=�Rڒx`{ã���xF�*���i�ReS���U�-�V
1�B�����-{:Ǖ5	���s�g/��lx�����C��,�H*O��P���6)��\�:�G�"�
���`d���i�7"�˨����a�S�f�vsN*�uЏ�*�T���1�wbӥ�Ĩx�t�����wȅ�n
B�U�P���Ln��'��3׻�i)��ް�R�Q_'����� CEj{WL��[ʧ�F,�o�$�t@6!V�VmGD�y��=µ5>�v$\�I��EᔧZ�#�ԧŜZkJzl�B�cL���5���=������:	)0@@ݗL����z�O���ɩx0��L��Y�6�lO
b�h���Z�mRwI��h@���8��A���kܴ�s��i�K����C"�8m�\o�ϖSL�A����QJm�,�4�1*c0�@c�qC�����8�fy�ֹ G������6Zʫ/��-Z�E�!��݁6�S�F.�<�l�<�"�#Ye	F�ٿ�g����|2z�%4S+Ҋ���	آY�;����<SHmJ�UJM�`xG�h>�R�1�^LeO:������Y��b�b������$SjI��Ւ�'k���pSh�cgV������d�Q�{U�C��3V�n�(�<����kHhf[���یR�iȀ��lT�$�3�EV����ʍ<�1���a�"�+�CU��8�,�9�f�?*�yۯ�\H���O�:Z�ξĒB��A�~!H�󜍪F�ߵmY�I�^dll=}�5�VdH��|0h��Etl#]it��da������ƽ.���v�������+�Ֆ���&��.�0�Ϫ�q�cM�H��s����c9=���m��r��;��j�2�U������^�]F{,�,� ����4�.Xo2��)I��z��Ō�Uf6�}{�@>Ec�Қ߱c��$�9$�����=�*܊X�Ji��)�������g43���z�u~�e��n~��K>8��A@{�ݱ[!���**Ԅ( .���T���A�.e� ��|���G	:#F7ǏEf�^�Mu�\�we����ù]��w����\�vqص�ԯM]1��Iӕ�CO2���1Na
�{N���@)��NG8;��:��*���{�u�"�GX'������D�).��i���Y���ZC�q]�r����|j�-׭O�A�� yd�h6�9�X����d� �_�X>�~�K���_(yE����~U�jCzj �Բ��oʌ�S<q�����4d�ʑ��[�A*�t��&����5�;s^���H��uo�����	��w���+h����:�E�;(8 �AfE�Y��2 ��7:������`l쇐4���J��Nbo���[P���UH?�k�I&$��'��)��5B*�[?
���.R�܁-��K:j`��(^=�m���)���$<�U{�^�fS,�x��V��tUb&i,�c�O.�`�eX��*�3�P�3�>Ֆ{��(��S���-�j{�U�dE�-k+���
T�7Q��T؄�N2%ܹk��
y.x�<aƙ�ɜ��B&��P.��^$.휢I��`6h�|�����bO��`B(]�I �~>y*�x�Y\� ��a7/����Z�v�T���[O����r3�$/�~�0v�sp1�Ũ@K��o��.P��Oր��y�6$�*�
5�������|2�MGڡH��r�y��3Ļ���}#)�P�9`.SoY���HזWu��R�-#I�2��aony��J����S^��b��kgh,�e<���Ɍm3! FP�i��or�B*۷b��I,�f�oF��J��^J� �	�{f�gB�Squ�]h.2@Dֶ����#W�Uߔ��=�5��SJR��ht�R��҂�4�'9A�{��$K,����/���JƤ����``ô1M7�dxn�YJ���/�hqu���a�\ip�ztr�Ȉ�Vߧ�9LT
����?���y�A�2�]·@�#��әW��j�w}��f�'U�6���A������[�n������B{�$lzt��> ��W�5f��nJ*�F���
f%@����jaT�����`�+x��bXpփ��FЪ�Rs�υJ_r��f,D�8E��C�w)���O,0�/l�jyV�"�.j����O�l��Q�<��C�Qrߍ�Ԟ`π�V�d��9�B\�^�}@�>FfC����I����Amd���'ѶB�3���T��MvKt��ao�	�Zq�h*���pN~s�P�i�&j�rls`&�b$���5�5����q�ɒ {7�6M�L~��*K���aL�i�mqh���M ֠�����l������U�|���*#�Q[p��?÷��:�K��\ǧ��/r�.����{�aFM�-�%7����ͧ��Xv�*�F��>���2�� 0��p�����)kȜ&�h|�o�	/Y�����w*�PaӐ���K�Q�Q���7��;x�� ͺ�����a. ��./�*�l*��n��ÍxA�e��^/� ��}�'!�[�?���7�d��� `x�fT-Jz�XO��"���J�d��F�c"^�],��{���}�e_;��#��hL�F�ζ�n�����妏f���nKl���l�ef��0��zE��!��)�k��AW*e��S4������ū�%�9r`���)��#0��ī�s��H�Fl�J���K]oX�}���T��5��Cן� G�ɞb���M��"n�"�z�S$��v��:�FI�5{���¤�]k�\1.m��ѓK3ŗ�*�O�ېѷ�:}1���1\�g�dn7gKR>��-b���,)q��PP��nTJ�� jݼ c�R<�&c�{"+r��k�c���;7#��i����]�m�6m��8N$�-��vk�щ�B�Y� T�x���C<�/i�/Kasg.��/�	'�SV��,ͽW~�@Ԋ�����*�qp�`����|ҁ�/ȘSp���`g��y��=P��b�l3|`��2�`3ǈ�q`)K�$ rh+�J`ZOo�L��BYI`�DH�n�(Z����	bވ��.��|;p|k������	��/]g*�N��!���Uءˆ���	�2?3���MAdD�{�[i�B{)gb���M;�/��E��5�_w܍c�����?(�7-+����K����Sb�:qX�l.2&��
�2�U�p��BK�&|I������A���*G�j��.�Az�������i���S�@c�`�R)I|�:zҭM˻>�dQw��o-ak�s��#�_n�L�������,��L<զa7�C��}[#�t��>�x2�Ԏ��~xO_������2�:�:ۮ�򪭅砖�p��P��������/�9ri�X]�>p��"t%M� �'r^�lN@4�����ϙ�"�K`�(I�iX�{�ZT�`Fxs*��`ĉ`9JⱧZ��nNg�B��iSJ)��ܣ�RݝI;@7�]zL�㊄�qQ'\�5Jn�hW��b��*>�5F�4Z�W���z�L��Cәo�'���$�!���f��wyӱYf^��l�|4c�gƲ5���ޣD��\>rD^6��Cpg|FwN�[����c����"���]��̵!���N?���E��DU���k�Gx8@
�5#p�L��)�H���7���䴲�O��_=�Į3���$N(�K)М���КsE��%w�,#P=ɬ���Z��N���2������'�.�u���#%3�q��F�t��
A�wȂ�'d���7���˄�%Co�O�7�S[3�Q�+�U�JA�>��z����23�]��K�J���<�2�U�j�6s*枑�ȑl��446^W�F�֛s��������ծ��{�<?�pS��Հ�3�f�l�0������� ��s��s`W�A���/iD*|Y��{$rV����y:���)!�|Fj�@o����>�,�f�IS��cVͫ�@޴�iY��,?Q�4�7���,/ ��I����c���vh�a^V�m���Ӭ�Dyu?�\�]$MN�`�.��: �MU�<k�A����q|�ب�R���w�X�B���t�$����'2�+��@�p�;���4��W6���f���r*j3�]_A�)�ͥ�^o,�D�I`Ɂ��6b�P�?q��E8S�|���GB��`�U(���ߛ9�	S��U�]��7������er'/ ��#��oS�C�%�@# Zb6��⫐���$�i;��~	�p����#�-�� �
®�-���5؎j$ERbϔ1w^������5S����\���`zt�����r�L�2�#-��&��$ew(�r�Ê�:�p�h��k�hv@ťdWa qC��C�����MH��.)���F�f�:�ފ�"%�B�%4�8Ax�vk�Jx�l%�M�f��N�8n�t��2�3�Ou��ML A���{������i2]G�5�_��1���iZ}����<c\���ow;Re῭d�bK߼.��Kk��!�L����^�z���:o���K�B�����/��Ջ<O�a?��/�VZݝI��h튔����\�w�ރT��3��W�B�? �Tt)LU��3��ӯ�0�)"�%Y|l�QE-���÷�2o�k)�z3F:hi��Och�emR���mq|m��iG_��!�Xo� �$�MΗ�ST���w3j��䜽���Ć��7��}�U��HU�U�sH�k��de�t<4��s:���։�HRIrxG�ֿߨ@��Hw�g�v��ɛ^܀���`�ĥQ��K�`A)�Oh ��ʚkd���Ү����w-
տ�#K[t<���x&P�6�!
�¿*��\Cg��9]�=ߕ�\��P�z�D�-^nz��.�k�Þ�{��7��5��!���z����ـ|ټ�D���F��k�R�1���zK�<ĺ H�����"U.��<y}�8�
��V~\��IAS��d�K���햒WC��צ��P�my���ۏ��Y?@Bp���,�?���N��^[�{h���B�� ���a�t&3W��k+��W��ϋ`7�?Q����;�{\���~]B�Zu�<c}Δ%��iE�e���,��]��|��5�����ijMt;_hmMsfI^]�u��T�ӧu�zĐU&i�vD0H6`��
����N����K�[��_�m�s��àT����-�0�6�7̖;~g�ΗP�� VQr�s���о�T�r��@ư��Ҏ{���K�w��<�Ua%���/%H�n���Cp�1و�A�6���XaFh�Mc������6�"A߁�z�`z)���#p��w�(X�?�����_Y��Z�JrF�`At�q������=~�3
��#��`8jsX�`CU�4V��8�WA�B]{Q�Q.��܈X���"����yE��t=K���b:0,��r��/��V�ftz9�dL�Z\��*�|a�oKI�U5	j�BV��$v6_�I�,u����b���p�Cg��%FgAlx��,�~����0,m Y��5#�\(���*%�GsT������y�5��& �z��k+Wj�{f$���A����7�А��~ u���I#�D�b�@�H O+�\dh���ZO��H Fp9P�}R�G��9jW�
��U770��?s�XAގ_��q�B�)����H8݅g��l�{���_ j@(���}�P��o�M��S��{\DP���x�;��0�@ 19�9~O�|�Vu������� �o}���;[�S��ylX�=�4L�a\|a"�����D���O� [�yk��,
�'|���ĂB��v�Q3A��X̃t�r>H�k�3��D�06�O��'L|2�ETYFm^x]�T]\�����cZK�CN��E�!���$	��w��B�Dߜ3��ٞ(G����]��s�\�d&�����2#a��M�Wp�n�f��B�kdf�M�x(�r)ޢ: 6?j1�~ٝ�z�HĄ��C�Wh�,Y�P�2�����4O�j9	ɰ��PIF�AG�++�C��1�V��������gc �
'(�˕���Ər`�	:8(���_NJ�x F�\�*xC����\C7��2�<��wM7�R&��\������ˌ=%h�R`�nl� ָ\�g�r���0��/-�Crρ��P��7�>D�:�۔I��P�Fȸb�e�潩�֓�X�D�B}��ؕ���e��VL��I���ʋBz�k�a_h�1����=<p��P�:tRe^	E]��x\oRJ����^�q�i
j��|��2��Y]�(��I�UE�x!K�7�=��um/����U��-��7��|΄l�� 2H�gvI?��k=�]̯��ׅx4UsJ��9b6фNJv�Z������6\���i�c��?�����2>=j�j�a�83ӭ��EA������#pJ'�!hn	����̇3�ˉ�V��2�O-�,ƽ�S]@��n0Y@�����\~Ͱ1S�~�� �w�?٢���F8��7�1��.�t{Y���4��9�M:ޔ���j1�VR�����͎� @8�R�I��s44��a�1�	6/���􇀹6������D��2�>���G�J�*�it�w2ׄ�r�`,�eؗE�H��BI ���� ��gI�rM�&�k<�V��N��y�����S@{��#3I�9����d�_���Bs&�:��+������OT��,������8]���y���kkvѦ���6�z����EK�Ss��/~�#y�����+�q�M�=�t�;���<��c\E�@��%w[� �.��C�|)�	޿���T�}'0�S�3@������4���o�rU�����iyqQ�j1b��,��5z��X����p���m�/����.mx�����C��^���\�K�Ծ��a^5J��)[���Y�E�H�DAn=�\�� ��Ch�5ۢ����t�L���ƍ�?��b�9rչ@] ���.L�7�	p�T��d�W��~v��4�*|��ZX�Q�*,�eD����o��q�t�v'�7(z_bh�����(T���NȻ�h��H����vÑ������0$���~l�@��:�ɫ��0`&�T|�-Q'КG�>Ee�_y����
��'�>�=������~s	h�5�JGc�_�MeH�`��t�-�]q�-��q$6B"�6䢊~���O�fmL��J��-CX���E��,��/�n�okl��(4d�tՎ��3��1К�#{7֌LL*
bA5hl�)C�jn�J��� �突sR\�K� �� 
ֲ�?�^_	��b�ۇ���'h�K#�a\��G���`Kr��^V��Ix�o��Fh+��wU{wy�f��8ҐQYf���M�]�ML2��eχoQ�G�j�p�����ѽNSc@�����Y#?	J�'y-O�Ka�\^�O�j�[(�lc���Re��:�n^c-֥��q�cqN��=����&l�ц ��$��ǩbV�>�.;禠X�2\��(&r/^T@z�l&w�[�Ş��x������Va.�EcY��i����BR�jX$a�n]����1�!wk�����A�(0)�1����L���`�8�' ��
�pp���ߴg��U�iP�	���ƚa^��,���SR1�g��g4��V�q�N�wk���u��0m����u
���4������-]BǏ�٨�3�)�N�WＢ�^��/l!?�D�xN���-�c�"�%~0����)Ӧ\��Q�������}�8[@��q���N\�&%�s�R8��.7����sN�r��zG�G��bj�mڬ-�g7�!���y���x#
C�-0��q������0�,Ȩy���-v_٨)\!�[�|F���8���=}���˥b<��Ʊ�t>���񎞷/�jp���NI{�s^e��gχ��~4�V�2Z��7����NW8m���b�ޝ��#��gWC;=��*v��CH<�2�wJ�l�)-�o�6�����;@�w���R����Vo�@c���7���Hp�d���R�s.S�>:eiY�z��q��=(�J�h�yZ�n�YL��i_þ㆗�md$��5|���&�2���� έ�GI�0�N�U����~ꤺy�l�X�8	x�\"�ƌ����Y��c9��ɞ��*�RCغ�T��ᅋH��(p庙�t��z�y����N�<�
�@sZ�\�,��f��2{=��ƣ��5�d�3�j��lq1�d�V���?�*�fK�-0�z��D�{����>IèS�&�~ߗǻ�h�=�� �ډ��~$:�Ÿv!~��+��6�d����q�(�2��k8a-߀�`ÞL}fw�۫:g�@-g����'J�=�?u�����U�'��ŉ�ވ�k����ߖ��H��ĮTd���#+��sdJ	~�[?m�'\%��đ�]_�1Ѳ�r��l�+�3+*�9o��o��Foco�t�V�D�f+;&�:����x8�H��]�d�����'$�M���f����3�FK(��Ũ��Ep����ֺ/�WmQZo�(�zsQ�\$��LO@`0@m%�����P��Cɧ���oACӞ����W�hJM5Vm�f�K���5�@����6^M��<�	'#a�k�����l��7�9yoOvz����OR���mvE_���.d62;���V~z�7���v�?E������>t��ʐ)�01�u.�������C|&�S��� �L+55�덌ἡ��@�e97�d^g�vp���$��iP��sأRt[0K�pCn����*oo6���X�쪻������vW�R�D�o�;˾����heJ"��,�����߯U��'T���q��=�rF�4/P%��a�xX�֖q�z���8�[&�qW[���O~�1����Ul!<I�g҉���XV�ǰ��}��0�|�.¦��{�}�*�S'p�gf�T3	�?l,�\�[Nl=��T��%���g�!b�������d���ۢh?�d�w�B���Q�!ǹ_�6	�)	�
:";k�(wf+Q~o�C9w�!��O\�O);�}�i�&H��� o8����=X����
�<6�i�1�7l	��`v���	���pK�}"{_�%�����L����o�LB�ฯ���eB���!|d�㥿�8�Y؍,�}9a9�\���b/h,J��,�o�%�6�����OW��1�r���n?��6#��\���Gx�����ٳ_��6��{y�U��A�����WU�1 ���0Ȝ����=@̺P;$�t=�PnҔv���LL�PJ��Λ�W�S5��5A��)x�d.�.6�e��=e�Kz,_�j�� �	X�qH30K�AL��ĕ��Tm\jҢ����8������G�(������akԇ��@Ѯ�ZZ4�]��T�V;�\�I�]ű1~r��x��P��������n���n���:	�����d\rM��~������ī�`ˏa?д9={T����
�};���ҫȏ�9�1�e�t�k����en����������s�t�m|B��tX�6�N��~W��/��8���QS�jm���ӷŷ���{��$��6��LQE��4�,��
<,��%\|���'�7�Զ9�-��Gm.�!�yf3��Pl�v��Ik�<I	�x�2[�:&9�iT�&^��e���`u��ݸ���D#.���H& Җߺ��\����ϒTsp�{�5P-��P�1~�i� ��r�d"l�/�-���}%i�e}ȵ�h4J���~�EI�Wn��A:S�;�P'|�	s�M��6���I= g�;H�h�T�ilv^]9&�*_Xx2lFF7�^�����6j���M|^<�.� Z��{ku-+�̍�3|^#���a�=�(�Եp�s���1�N)9��.
�[n��{G��DY�ܜ
y��jc��*g�,=�nS���l��� y�)s�̞-t,��
��k7o׻⎾ǩҁ�X7E�	z�#�0A;o+*$�AIt���g&Յ3k��|tNG���m*�����2Ա6�eN�wt��y������4��.�r_���A������o�D7�)����I�<�XR )P(�prAǫ�((Īua�����j8Igp�k�d�z�~Z��Ѹ343�HI��C���y&��<�~F�]����{�ױ`;K@�/+�m��@���E�!�q-�1��������ص`����$|��o����G��ι.�����	��:fy��`��>�T=����������pxq�����dk��7<ym�5�� ����v}*�	��ˣѓfk56���n�^�y�g�W�ٺ�zMؿy6/OiT���M৐�5�j�-���ܒ?}h硚���0��I�����L���!q hOZ����0�W�(jƔx�KkQƎf���ܙm��`�}j���J��:+�R�ₒ:a��^i��m��|k�_�r���� d]Q����)�VE��H[�/�	���:���K-*g=q ��İ2)��d��>?XцWNI���a^����#E�D���5<,7>%�~&���%�G��bs�@$>
Z�x����!�P�0���K?S�+�;߷���!Ң�o���MOWʲQ�h��H�PGTj��b�L�|��|�#�K_rwE"�}��������'<@��AX�E�/�MI�mA���v����*����$Hu�Q�Od����ݙ��X's�Qwԁ��E\I�X�R�x�a��1�qJS)5tA�܇�H���������1*� ��uY��}�`<��#V��)��f"�z���5$�c�̄�hL?ظ9
s�����2��L�g�*Pi�MXێǚe���*�bnpP�����-���[s��G��b9����L���a��/���~mAeb	pMh>^Oh&�3��X\U'���e��*�˒
��/�KTc��X�-D�VP��t�>H�MypT΂��K{��[�>��^�]����TM���؀:᧤�jx����*&Ь�a���L5^�+��w��Sm1��iF��ي���x��ݗ�T��z�9bP�N阍���3��p3��Q��>��E�a�w�<V]���3��TX�V��4֓���e'ze�Y�b�~��li�$��-HU�(��`88�!�>~��}��'0!��9m��	xOU�@�K�4��wu���z[s���@_�T5�H��ŲQ`\KA�����jJ=��5cD��(5j��l����X1r���o��?��1��@d����$ŧ1=i�/�����O�2-i��\�o!3����SOpo���үp��	���tz�[;r���E����p���t���E�ޮ������C�����G����<Q��6t~Q�0�mV�K���0�% FR��ӹ��E# ����_��&�Đ�nn@>�.�
��ME��3��ràF'4H5ց$�fF�{��2�.CŌ=��2�kP"ʫ��|��Yi6�[�r�*���˩Dۊ@�����v�.}'c�v�Y'�F����� P��*t�b���G��@�.�%���C��\ю�g�ƃ��%�"Ɯc��n�x���cKV
�RzȰ#�
�"?���#7�l  ��*�
��C�
��"1R�CF��Jr���XT�O���B�#0�ʥ$�&����s��N��`�F����%Q#ނ��=@��maխ���E���*���+��a��L����F�kK�����S�T�
R��7��k�Ͼ;�n��3�*5��Z�
�f�;�cYw��ݲ+�^M�?ך	*�rkv4,���͢���\�5<9/�xQ��������<6=�A)�<~�,Ӈ
Q8��'��kSJo���	�7X���O���� ���a���H�O�%|"�C/��<��ZN�h�>4���6V%�b=�	��S����V��,���8Nl�
�S���_B1�ت�A�s^zek������7,��.�S��K�ΟlϹd�m�$�w,��4z���M>�ҥW�j�M$�
4��y�]�W;˶�.~'�'4YQb[,��aj����n�G�2�",U��YF�(����$qA/��N�����D!Y�%Q3\��00����C��"�� �a������IH�ޡ����F��%/��Y�����
�n΃>&Z2��n!�-�۾Ed�Q%ZH%�C�Y̌m:�ߗ�3���n�k�G��Dz7�����#�����Zd�/��IGtH�뷷r�Ii��� ��%��;S��f㛣�����O��cg����;�.����!�Y
P�n�-�m�T��QN"���>5�B�6�!y  #���l(��C�k]�|%9px��2 �N�Z�X4q��d�<{3�{S���������/��e5*1s��wS�A����(�V�&��>o�Hh��@�fT��/���e[�����k�K�
��B�kM�8�0���l�TVW�+�D��[��a���e�G��[�%$Τ`����)�x��͘N�r���@� �1F��Kh� ���fD�V~1@�w��KoRe[$�!�[���n*�>�[�Y����2w��8<�2�v�`6�pE�����^.Z�d[��r����n��H̋��_#���y�Ky���ʧ=#��ܧ9���'���EY�#.�jDts��5��+�c\����rfE�e��;�-z����>t�����j�IA�0'��0������	+���*�]M֡���$t�8�^�r�)q�bJ&�C
6�޴h�	�WA��ϵ^WӖ�Þ��(��Y�rؾ��Sl����#}�|J�3u@�}��QѴ|�`���s\)��Δ��*}?��ߚ8�A�"1|�V�z�b7}�c V�{�Y�����f/�ݗ'�ǲ�m��He
@��x�c��;t�Hﴞ~5WZ�_b��86�~W��W�u�v0�`&�#'9M�:�|9����&�,�-Ws�W������y�|��B'��0��n~"8톴;�;���ƿ�������G1Ǿ�bT��C"�VV��د�B�z5��F5�y贂��I ���M����mRcOc���]�;�+.m����$�D�����돞R���E���a<[x���x�G���^q}l�wĘ��S`7������[�L:�;�������}d`jpȸ��QT{�PP��1��J�
�[X��g˾��w�0n���M����v�a]@�������:�Y����/�%�����׿hzT�X�<�k����+&��1��²/��[z�q�d}z�:Á����?YU���ak�:L�w����'�`�Z�3.�AY��d���U��O6`h����U����"M/&,ԫ1Až{���U��������ɐ�WS�ч����Y�ʹ[�;H�h�q`�Z�~;�4��<Ȼ�R��|f��Ղ�L�_(���S4HJǸ߲n���zG�ip�ʖ9�8
�H�{Z��*�Tp�ύZ�e��Pw�:��Ŋ�J��v<Tm��W=f�|�R�� �k@��(�^/�4���ع	�U;���@_����+�3cBUc�H���� �$�r��Y�i���Q`J��.�W� �CK1�(�i�T�t�o�{��ѳ��]�:Rz��ZȌ���Ͱ�����*�2���c4<L�vqt�V�H��2�'�ro�����0����M8�«��p��oE3D@"�H���(jĉ���N�E/�/w������|dW�ֆ2;�Z�4��F,��G�bs��Ly*�芅Dq+�*N�PE�{����[��=�r�=.����8tH����m��͏4�����f&5��> X���+k��H;hb�&�ym��Fy�Ʃ��h
�j|�Q`����BA��t�E����u�x��9Y�k+Df�����Gm- ��ٻx!c�9�� �߷,k����Ʈ/aVͲ��-�~�$;���u�:��2!r��vFb��[�`>����6o[�Q���W�rrg�[3�\÷�].�>G�1l�z��ƈ�b�Ne�3Ü�ya����g����c.�|������Ɩ�.��2�k��*%��t������?	���^�9(f�<M<�8�T�C�yI�4)-,Ό�l���������C1�4���8�;<������	_ԗ��+ohT���sDYTrƒY�[�p?���t�����|���d���P ��C�T�=������UԂ>!���eA9���x{�ܚ�v�k�&�6�.	 �K`8|<�K�sD�_R���W`�Z����ra�����l=�� ���f;�a������>�JZ3�29Wُ�ܼX>����{B~�{�O-یD,b"H��0LYnw��u|��Tg�m� :�%8��-�>lyU��-�������@V�0=�U��E�Hc��ʿve�ՠ����ģ���)ữ0l8�
�H-~,�	^�>��Q�����QD7����V�Y��1|L�d���iD�G�d�1�[�����؉�+���h�Cjb��o�r{��ɾ[���;[~���~� H1����J�C���!p09�$��1 0܈�LzbM{��^PG���D��z����H�A[��6��F{Iݶ�a�G��p@�L[�p���
���7�w�+�Bv�����ճB�ӻ�K��o�K-���o����٘f���B�~�}J��i9=���2-�F���u80��ҫ�8^��"B�U6�\.q���w���{L�%W�DC�4���ٔ�8zu�(*�� ��5��ݘ��%��N�A��P4���C.�����ɿv��a���25[Mk�B��#iIf`23*�eif.���=����A���9�8��o�D��3����D�	��?�������������"�lH5�³b���	��Q�N#�u��ѷ�_���lٖ0�N��'_
,���
꺚z�y��LJZ��w�i��ٷ�JfNTR��rM��I�����2ň�� h.+Q���r�t�V�h~i��b�V�nĉ+���t8�Od��J��-ٙ���B����V�#�^faT:���Ý�4E�=�͢�����0"�17��$�"i^|��mF;����z���A�ǵ�Č��?�lxk��mp%w*�AЭ��vODb�ֻV�$��Q�ҫ������i<�N߹v4���#5 ���w�p�m�@�_-��+~4"�5�kP����@'�u���7�>S�?�·���2��:�������@n�_F�	:�b��T��%HG��SWHG��R����l�PZ������-
��3(���Ϊ�?��d(��b�X?z�3��buG�u�W)K���fH�=b���;��_IH����0�5K;V��?A2M�j��]p�Oܪ9�5v&T�c�J���,	�A]���k��po���U�pTˮ_�=ᵒmE����j�J6�
���p�	Xc`;딩��e`�q˸�?����Q�;Vgȫ�ƨ"���ٵ=��4F$�o���i��2^�A>Ǎ?!��4�f���|� d�C= +�WJ����d��TRHg����/��)�l�w)��ȝ֬�k�D�8*�!m�8��|.<q�I:��8�,���EPb���j۞D�"�=�AYn9(
Y�ҋ��ob�nr'���V�N�ơ�Q�(�L�D Q�)�$Pri����IR�H��z�8��F��Q^2�,=?�q/�s��
k�������tt��H��DTO%֧
Q��[^\}2�0�u�����}T���>��xo�ਠ�C>�]R�#��d�����'ˊ&e��F�~A��t^1Rvhݤ�㻓mב�):�>��%�t*�[>��IA�&��wX�~
|�'S�1;���H�����F�=%�r�&;s4&���چ������̤���q[h
P��B`�P BX�\P��cD]j|T+��v�Mv��`�V,��@	}���,q4�C�<�C@�s|E4A�iz��l-<H�8B����~L6 /��Gl(ҶX�e��D\�뜨7Gt�}0R���v?�҆���n����'�=6�B&�-��Z|	�@�R�K\O�>�D��&:5�������q�@��DE�X_�4�� +���m�o�G����uy&������	����#���6ߺ��!p�A!֍��͈$�c���;eڍJ�S��(S,OB�Ie����� ���PoQ�pZ;Cqh��a��M���w1��&�����7���Ǚ帧뚅���gZzƂ��߾ے�&p:I_5�䳩MV��+��h�s�4�d���4��K�z%؎b�z�M��<I�(�Ԇ�����P̈P'�G�ő��,�9I�63���6Q�WV�H��T��^�`�g�Y\����~����)Q�\9 �3~B4���2w	�����3B�x���qՅ@�;Ӝ"s�Ӭ�P�	]��n�l�9�=HAn�v��ĺ���h�Q��#�.�h��P�a�����m��S��b8{&%�B�r{��+�꟪�=yݔ?�ղ������2������Oo�w�c`Z���V�_]ˉY���_�㸂C:�z@�pſE��P�M��7�>���0���B�&�_�d�hpW7���G� xtzz�r�D����$)oI���ݕA��([�g$��J͘pW£�zʊM��6�x�j*�`�5=�k�OW��k�9�T�o����x�/<��aU�T_v�ۥ�N�qj�Z��ŝ�-2��D��O�1#�<Bˮ��(���5i�d!jǺט�Qқ��RĶa�>��B '4�ߎ�.�;�+���;��b��te=�y���
غ��%��[���_Hj_ǲ�Н��士��\5I�QX]�D~�7��,td(*X�d���aU���(	?E���q\
��/O� �}!��3;�+����������%I�%���4����ЋHD�7�s8�����,2֜��p9b(a#%";�ذ�A��;�m��P0.�ujC���9N��38
g�ޚ?�Qia_��!K��m�����j�}�� �?%�ܢ���7�R�]C��Ŏ���d|#����&�s[R���pLs>d���1�}n$8-�{���,�Y���tP��Bef.���8"�z�K��Ó&Bo�%��,�,��AsK��_�(�u��
�@>���O����j"w0��,�:�י0o��)�<9r'�b�@�* PҶ�>��N�bf=J,�C��n�~�� ��u���"�px걅BE���{ ����xAx�w�4���]�\�xgU6�F��89�N������C?���8�i�fK8���E�&��@	t���^2.Y��:�����Q(�)E�/�\o�������۱��8Z!�d!%�@�|�/�a.牳5
M�驙1w���F�������WP�/�R�C�̋df�I�3n���5Q������**l7����b�!/��q�,o�A������n
���ܵI��';߸<�KE�N��'�2�Ty| `���A`�9K@E�9f��I*Z=QR��)��GQm ��,H�ǓF$��XѲ�˶-�|W��iYC
�S�"�E|����]7Z���b�O]n@S�1�ˤ�֔������"Xٖ3���iDAY�~h<uhj;B�e�(L���M��p���TO�y�����,�]�0Q6�gf�vS9������TH���U�Ya�����]{�?�^��#�m�����`�z;2���0K�͉��WN��M{���}k$�����_є�n�u&̌)J�Ѱrw:!q��H���Y<Y�}�p��y��Ϧ�ߧ1��bH��F[{J��w���!/m�g�����Φ��v�*�����*֫�e\G8o���쓖���C��n��m_2��es���Y�pՋ�X:�����Xj�!7o��x$�V$>�=�z�����q����^,��I)!lȜb2�*�������"1�F�P'y���~����F�����'�WH�+_�"�;���Q#��F0�\�s�h���l/�O-ƿ�E��dmv <>,��Qm�/�o�&��-Z<��,���^&�ߘ2��`逸��,�f�'݌s�
&pƵO�����o+���/-�uc:�!�ܽ�^� �O�[�_�G��-	x8����R
R����IոbY|@�@�l.X	)wM�-�x�^�]Vܔ��c	�D=C�"�]��^��]r����p\�(t5+�1v�V��O��*Ft*V�E3\a���<�߄����-�u$4�����v��n������ ��?ޗ%<�w�~��'�z�*�<��䞩��1� 0�[F�Ɏ+R;�L�g�% ?r;hxm�g��~�"W��Q3�8kµ�L�O�Ӥ�/���a�=��+�(������Sqw1t�b������z�ˁ���?����
g��7��H���R��Y4���'jP�Ԝ�������?������; � �"�2y�J�z�m�#u��3MI�p{����s���D�Ȥ��3�5.��ooy,5<99@x`�L�Z(gK�<5uQ �/y^8��M��x�z��+8R]8���,J���'Xv�>�O��L�����!�/v�n� =��0��۴���S)��HdM����q_7���Di�:�;@���[MУ��-1�Y�]j5�R59 :%2
�y�Շ���Z�9،�}��&�գ�8�)�@T��%!���r���/"��PX�LbvRW<���9u���H{��;Z���X-�V�H{�	 � �'�ٶ�h�}B�2�k�~H�F1�4@}j�F�6��y�dD��c&�g{H��;@'[%�%�Kzk��{���p� ��7n�[x~KV�-pl��׾HS{e��l�"�+łSS��������U5�Q��ɹ����>$^$&��oqs0ڝ{����,>�A�4'S��ڋ�]�OF{��R8�8X(���{��^��ak�>�tL���+R1�ߐ�|P�I�.��yQ��=�2��k?��́"��W��k��9��#~E���L̔�|.�}���~� U�������j����e4ř~��g!s�@���T`i��ԓI����6�t��b�w���R��rT�"U��T��pS>������+�����r��}Yzg���e��@-Yd��x���ȏp�a|a�N�ct�?��C:|����n�k�����������3>��b1��,7���\gh;�%�H��"RC�9�"�\��P3�\A�F�-D�P�� r���?�Z���\Uu��bV��7��X��89���f���J�P��zf����@ �U'�mP3KgV1m�W�J:�
�-	�pˮPZA��<@t4��;5�>�MR����W���X"��Pq���Oc��%�=�2�5@�ĠrL�k��*\����9��>BG��D��@�l�����2e�ʞ���*H4��%m�K�;�:C5�{�(�8dT�?����g=�tc>���!�a�D�F�.�X'����Q��8s��7YWN���t�J��ͯ��߯p���P^|$ѿ;�w�n�t�{��,��
΅� /��2�l2/���'4�n��eѓ� 3@�EθE$/*��h}\;lu��ȕ���DN�>V���"c �.�͔�q�d%�V�s#���4,�L%m{�F� 9aS"���w&��[��1/k%��d:����K4Ci�ֹ�#���Tj̊VuC�Q1�*�+���u_�� ��ֱ�Է�����V���F�aSpԗ}��)���|l_
s��V'�3�r����P�.S��6�qQ��ab,V���s-�l��N��Lu�y�/y�E��i-�UD��EK�"0�\rBq�u_��]�ǖڛmf�Va���,��4���8BD+�l%����&��aNO�D����߀1S$S�\�4Au��	��+���
�$9/����}{-rx�C��r��e|f'���*��}��b�1p�7�I�����2��A��A(��y�r����sw7_�f�XrT]�I�xR��!��@�������B���,�P�����^�'�~��V��������/�c��`�~L^愠��f����I��t9��	�"��/��@s��yf�ߙz���fJ�y�mV�QH��U�7�g?,��`���e�cd�iR،���y�ݓ��+�����h�,/%���UJ3��C�%6*�w��%����\��RBƪH�^�Y�|�!}�\�<�bvvw9Q^|�̐mٱ�5�X��|,ݔ�zC�6<ta؍����R��x���[^�RL���s�<:֗e�A wb>X�E��!&�%�q�,�E{�o�g������<� ��s�.��N��q5�wAcC�b��}��
V�Ci��7>d����!�[��bN �M�O��=�X��s�L+��Od��oM��6�0�o�)�_�yv=L����-�d�`jα�'���������8&Fk�SH���*6�,٩FP`L+U
o�c�t[܄
��<���e
�\r�d{%>9�h�[1���]�u<k�&���`>���Yl�W��*J��.E�]<��ݮ��Y��2h+��I��ՙ���<o�6����N��]�=������_dr%+UA���\lň��ـ}�`\�g��i'��fd[�� r�<ͧ� ~�p��NO$�\x�uh	J�<������˓em���<��5g�9��3���+�q�ڮ$�p������d��Nc�"謍�U�b֜���q�.���.CT#��c���%�0�f
���Ǧvz�⑐���C32�O���K  Va�Y��CCJ�)�'�Bi'!W�G���%5R�I��ӓ܏ "��آ�P�]�w�<�Խ�V�ԣ�3|��ZI	;����'r�B��lPzޑ����K��S8ܯ��M�zdK�\��r���]��1���,��$�V�P�P�* ڿ�9�;��Y���؀�X:8W�`[0Y�Ӷ�bo�_��U�t�{��1b8����RX�A�7�t��bAJ�'~\n)?)L�w$y\�m�$�ۉS��������=�K��&=.�Ǹ�T)�&ږ~N�k���O|2瑑E���{V6��,+��6]i�ݦ��Բ}R�Ӕ�sYKGo��C��)��{��Y����P��^�t��h[U_�_�M��m@��"���'%A,t���h0��a�ĔN�!S���@�0�ꊧ6� 2X����)N��{d��^� L� Ues�&�j�y�>�"��a��+>E�^�͞�����c�ϼ$�P��2���[����T��Ü�U0iICz�1�,|���'j03�]`Ь�E�2(nh2ښ��o[���=X{6����GB�z�\�T�q�q��z����2���4��a,X%s���_����گ3��>�)������>ؚ%P�74@Nn����U��Г[�������������ٯ��"�K�PaIû{%�Γ�_����n$���Ho�Y��;�ݿCՙ9�U_T1,a��;S���6��}�$zA�뽈' �(�'�Bq9�_0�-fDH ��|t�*%�����Jpk�s#(Ӿ�����A��y'�&/&wę���:M����n���6c>Y
�r��F3�;�[^/�Bg���њ_�[+F6���8u,��\eK[�᠀��?9 $�8߿{kR�:KZ�(�}J?� r�`�S��9D�Qة�ʥ�\0H�<I���Ы��lu͛��z}2L�Q�?��j���=�g��M3Cnsu�,"�%_<�(�~�
���A<��K�ԝ:����Nv�%����dsZ��&:@��x�KتW�Aʹ�2���Ѩ��<>�	v%�Dߪ%�Z�+!�9��z$#�Q�v ��=���,,C�w$K�4/�/V���������Ns����P x�gל���^r5�@���J{d��af���V��20�& �AҔ�\|�nw,8���d�)g��􋕍<F��v�_I��	"�Q�,����f����\��L�b�SW��q�v��y�mhi�m����ɇ�*�����O�����.�Ia���v`������J�S!��Ԗd�+'ek�m�U����k��������ݖ���j��Գ�>FM���:y�v̈X.��?"o[m	��|�p��<����6�w�zΩb�h�y�>�h���u���a�u�i�����x�0Ҧ+埻��|��_���b@~�<���>�cA��s��Hd����*�tb�� FJl�x���wK�7��6B�7��}�b��|�==�~�?��*���h��Z@H�Y����Í9��s>�4$���M�ꀽ�<�D�2z���}�[@��a��OI�UKw�N�: �t+�Ɖ�y5��MO� Y�ӏ����+��cf������D�M|�I;�(.����I�G`t�s�po*>)"X�]�!�L��2��)Bl�&�ϫCV�/ԠE�����	�	~�
=��������NJ |�a��+�t�f�����)M�%���� L�X`pǽ1��΢�"l6���c�Z�����T<�G�ɺZ!�!ᆵ���S�E緟�'��):�����B���g�ŷK��fL� GV�4�FE.i���?��y`����4HHH�3� }�ًadOC�By���l5^{`$�+Og�剂d�-E[�L���sh^��[> �ƕ�Cl@����+(ɷ<VF~��c�okZHj8�����p��:�.��%_�@�%�ѠZh�+�.�1N�(U���������qP���;)j��N=�U���-P�GjQ�U����°��ܭ�)����Y	ͮ-�[��S�$��H�0�w�Y2�����z���j�q�{D�ӦP�C^�z�z2\F�1_/�iZZ�`p��+7EV�i�g�\��G^M���h�`�G�N���6��!F���lq�0���(���j�x��fG֭��e�X�^L��iMY5��o�C_6s1J�v��Gk +t�� *�	L�la�d%ن!W�?o\aە;T
�~�D's���X�K�H�)Z#az������{'�c����'��H���u�gc���+)݄�����[���a.��G��@!fHӟ��C�XTxy	�G��R-l��f����X��y�oN�r2^�J>��wr���vXs�9����q�[/¼���A���2�=<���Fذ?��"/���vL��Y�}�y�$-�(�)�s-�{*�m�}`�;M�ݤ=��zD�ˠ��i�9��qn#�ݞ�t(��Ƨ����s���PD��?���=��%��3�K�i������a�d�/D��.�e��kY�[�B6�����7���,�����tulb�|R�:_��{�>�Hi�4���~̹]eh���^E����`n��X&pc�����f��j�b�O�����Qы^�Zv⿢��7��'
!B�V�og]����.�Tvy�.��x8MN���64+!=u"�RR�5�pP�j�P��?zY�߿-|=~�>u��*��-�/�lv4!�<��^TO�t&O�v�7y���m�!�"/g�
j��!=����ﯞ��^��DP�EMd�!j�	N+q��)-Į�~cɲ�N�q�㔄3�O4���B���e��y���'Т䗵��0���|�~���O.gˇ��5}ؑ�C���
3~�4:t�XD�D��!s��=�f��R.Φ�GJ�I����=�^ш��TZSu�l)=F�G�,��d�C`�`Mc큁��}
�e��ss�71��:�����x��nC�
��s����;�d�Dh:�j0�������P�{�:���9E\U�H<>�ɑ��,�)���G���_c5���-�2)�v?��H�_ �	����A���X:z�a_<���E��{�.��Z�|��8������B���.����Ukt���G�H��JFGPS�|�?J�h���e���)��v��W3e!�r���u�Ʉ�����pd���m�<�r�M�[%�N���[�� ڸ5�4����1U�o�0P_��j�"D�5�K�#����yà'Q�v���}�&�,�m��zf���q�x`_��.#B�m����
�)�ZN�d)5_UMY����
v��*��_�4�@ɭ�R��|��v~l)�ym�;������mkN`���RĞT�������T�>�Y�z�S� S��a
A��I$I䨁��W<���*�im�g�pW�'����p=���3��1	X���R;_Ir�P�ջ����I��l��xĐ�k�D�·~m?6��+����(z�n\Wc��4���C�*�eG��A\%�w>f��;�R,UO�h�WEg�}��d�K��{Ĕ#��!�u�ﻬ��]Eq�&?�C�]�I�~�=+�����hE�Ƃ�=�����\��+�9z�=�������P�A�Ε���V�6��h����`��W����a��ܰ����>�#2I��L&� w�H�*4��ԃ,|�$g'�6[��܎=�Gz�+V�x�/\2���$��o�{B�lw�dN�� ���G�x�2bۃ�t�$,1?���ԫ,�|�G�N'Wab�`m���r3��G�]�T��u�&�[���mH�9.�KB���]�aa������M�#�0�w~ɬQ��x����
��CFbU��n�����7wU*xS:_��/E5�������r�q��V�����N�$xKV�L�b"���E9~�g��P���Ӆ9��DE��&x��Vz�oU��*����C��?R!����� NHU{o;�N��uډx�� ��嬅�V�f�D�[+$��؃9c[��{F���L�I���q�N�U�'RX�C�7����M��[}=��ܱ}CI�������Vâ���c�,)3@���I�c��sL	�u̍,!�.L��,�(˒�*�-jm��	cqc?ۅm�hmR	��k�p��&�pgl�`8ؼ8�}��f��Y��<�1>�VK�(^{�m11��7�ϑVKУ�ka��������\��8�b$��e+�A�hWX���G���~my�8i%�ED?��TQ|�%Q1�w���)�4N
D��2)��o�����o�9��xzgz<)�wj�#Bvn�6�2c���Sw@-x�T�h�e���6���з�UvѼ)�>���h]p1�LRw�i@��� ���u�>�ElB�j=.�?��`h�g�5.��$c�d��*eu��~:�8��)G�o�c��7:�͓�f��s�n���P�T��^uA���RN�;(��F�'W�f���43u��H��3jJ
'K�KR����2�{z��Ļ��/-�@�����҂��2QfJ����v�I���]��X�%��&NL�.��\��n��tNR�8(C2)좤�DCR��x2TQ���;
kFsoR9+n!���v�����W�Zs��0]��Bd���3A�x���/���<�74r��.ȴ�gB�h�a��s�r}��xx
�Pm��k�& )��0��4W�&�q�^Gb�w�O؟|#SPFY(AL0��A���1}��]&}��,$!�1�������Z�5�8��ٗ=���A�T��a�J%�lg�o�:�c�Bg�l��O��|b�`yQXF��QĊ#gl�"T�<��I��]��,ҍ������X��V����z��Nm��lc��|��G���f�g�j���Ά#.��'�7���0�ٝ�+L����A��GI3�VHI����|�TE{���rˠ�f~����:>��5@b�*u�)g�;[p�ݠ9�3����F�x֤��>]r�?1 �	��/��D�+kXdb�>`mq빻�O��G#+%�(��M��_7��Oo/�󫻄7lL�j) �l$�}�ʆ�/���tHO�3Ó���'<� �^�\��Ô�m� ���h�T�ɍ"�t4C;�����@�=��b���l�~�;w ���A�=@2����V�8g�#K�sN#��9�@��i��U����U�e�� 9O�JtnK �3����LЏh��B��_k,�CS���@��mB�[�F4�K�U�5���'��o����y�.�L�dm-�D*6`�Nm���
	�߇�e��dt��j�J*�D;y�ڊU���n��Df1�ik��|���"*&0��CB�-d�`�X�~�S
U(X����f����\xM�uW���b���#,�$�!��֍�Q�RI�hb�����?��c��� ���*�S��r�H�&T|	4��z��D�c��@�ُsTc�.�����*�'�R���;���]t� �ߢ��mG�b��-�.�#m�&��={�L�h�. T�<�唜;��=�A�F�WHc��H�p�/0�!��U���2�X���vAG��Ê(�qkb�$���!{\���(9؏Z����.��'*B�Z#_�`��������V�ݾB�T����bx��1�U��I��ut%�K�nJz�����(Ix��/g�5ǈ�3��қ��;�up��3�Z�����Y�?u��������e�r�.�p�R��j�R��X1���w��&�PA�mC�l��(�����h��{�����ޙrޯU[/1UT�x��"�[5���6�e��;$u�9��i�O�����+@�m�+���tYm}�_u�>�L�ތj氃XX9y�)�	��a��"j#��)��c�;�`�xA^qRG��ײ�0����611`mc⬲�6����Mt��!�h4��b/G�?GUĂn�d�����\�@4 ��p��*��w;;^h�Ǡ옟\��N�O7��k"ޛ6��1�Pwé�D���7o����V:Ow!�0B� e��Ե)VPK4�]]���J�B�(sc�G�A���X�t[;{�T���ZlR����ˏӌ�y���o&��s��ɝ;.�N��$%�\��h��5M����j��}z���^#����Z����|�?�'Z\��c�\�xW6�־WF�j���E��j�Z�6i���?,3\���y�gD+�,����s�U9g�F�)�D
��ۼ)UY�Fi�cP��"�,�Ԡ��YEDɭB�s&Ѭϰ��!�����D. +5�Ye��+���l|���+�׎��#�)��!�B��E.牻�3浀�	}j��E����R�?�<�c�p���F��7Gfj�u;閳�"2��df���B��,o���_]2�4��:hu�����y���u/������ĨŎM�l�?=/���C�c-E�y��tĠ����_�ݭg 6?��0�Ni��΢lƈ*�������K�f	xy���`�1���7���n�^���T}j+|�g
��ܶ!�	�Sa۾�#!���i��y3jp6���QNឳk��s�`�� "X�A��� �Y��}��};Y�2�y�B<�x?��~��XI%ς�����|b�����,w(���uGd��aL� [�~��C�3�wǼ���+�D���?b�8���Y��Y]#���|Ɓ~��_�:����{ܭ��N����K��~�^��P�D��V���X���x���v4^"�s�k�1��ܰ+��+��vW�]�w4���XBay]2�m�u.��m"H�n��Uocِp�3�(ά����N��e��a`�_�RF�&�B��c�ssA�"���ȯ¯)�q���G�KGf���l
�������SU^�����A���-�
��-M��ldh�@�Ek����H�?2�7��1s$��j��Da����O��(�6O*��ŕ�!���@т��t�蔪r9�!{|!��G��ʵ>&P�_��4�	b
�TWZ)��xMɔ"��d5F�.�Z(p@+n�q��8����`�BE��M*�o�:Y2K�W�n�����ϙ��?�H�7�m7\�D��e��\<�|Y�DOZ;��z���-�8��e��_4��މ�\�9�G2ssj�{4�]Ю�	�0d�5w~��_ A�C|��r�<g��~���$��2����iq���CHؠO����I��#�E��!#��l{͜E�-��{�\cV;Z�(�!�e��K�&^20c���CY)/������O������LmTĺ��n�v�X�P���\79k(��!�lx����E���N�.M���p�ߧ���YS�\hh8�icR����H��bT�yN&Yp��,����~x9�YH�	sSr0��FV�ۄ�i���6��8y)��N��<Ϯ{[��#=���|�J���q�'�l�x폂�L�
���C�$���8�g"�;�`ǔx���g����r�骺���L}Y�(T���7�����m�AW
:ws����G������Nڒ�m	�Y�42�
���Xc�f�;�|6����~|�#Q�VHF]��j�8�,
E��Sfg`�=Zax8z!
������C|��}�~��t7�S(��Ġ����v��
�F��KR�'帟_�u97U�!��P�QN0���^W�6C�������Zt�k/[�ݑ���jC)�E��l��!�N��*�`ʰw F�w��7VWS�!�9��s�xE�W泝���h��^��T:�+r�����H����VEކv�BU<�eJa�K��Q�e���_���U�Cڍ&�K�N��ؠ��s 4�/�"��)~V[4�t0�z(�.'.�`���i�c��q���~�W\x��T�����H������U_��`p��^c䒚I�x�	WS֧�8}y��hG؋�g��
�'�*j�^��)\��~&By�YE����'i���U��W�0�9��.v��^���p�#�K�r��pE.����鹴���.�[��B��}$+�-g=��)��䙙#���GЪ�L}(Ș�GҷCL�Y��ۋ1�+�"�<=����u��К#*�D*��s���<t%�1L�>����	�.$x�ċ���R�GN^k���v_����鲻?�iPw ��4{a��R�76Q�숒���E��$m �bz�ot�`�s�uB�<�[:�D��ɕa����'� ���C!��39�!��tx���ih����|n�5J�X����#gb|"��Z�L�@�ε���q���͈��6�W��WN��(𵞲��<�A��GI;�Y�D���˪b�"VZ{'�+Q�I�?#� �U��]<t�6�F lCB@�Ȏ�bA�PK~-�����Hn�\;aP�^�w9�Y+�=��Zffv�OP0�2�?����tk��%m�ݬ`��E᝾2�� R��E�*43ľo-���C�U =�>�gB����EV��4��5���+�:!v�M�z��E !'�#�K��^�'<��o���>ъ��h3�C�w���z��I�P�Yi�\Y�B��r?�:0���o����q�$bd.�W����Qj���n����S�G�4<\Zj<:U��jH���lKx@�)����D�Z�;p�������j\p�\y�����8��^��O����C�OUЗ�G�	�)���>�Q����h�+;��/\������48��{}�R��F��;4�f��7�TN7G�@���h���!i��r:�(AE#1�������)g�'��a�~��\p�ΆS�����Y���|..Z������PA�`��l���g�=y�3��9�2�a��ק*����Y����rҭQ���S	XX���sACS���}���4_�)u|+��5����o�:�-�$z��"�Ʀp�$s�[D=O��[s%
�T�$*B�����6��d��N\F��v7����u��4����w�%�l��_OI�*����'&y��Q�&�����ܤzS���i�NK���]�{� �4~\*c ���0�]��%>LXu2ˢ �F�=hT�{?��rC�1E�Ι�9��%�Q�GX�]d<~� �V<�H�8�5�Q�D��\Ѵ}�D.�Se
�k�b�1� .�*�?���a �HX���B���f�Ky����ж�5��=��N<�eӟ����	+'��ԭ{��������"3��w`I�X��@�k�:��>�cLiA���6��g��xDz�P�r��6:n��( ���v�|����t���b8�z��s�z� J�� ��[ȉ+��Z�jNO�eg��Y��:��@.L(�H�xt)�>\V�W)�̼n�����2�=N��.˘}�����^3Z�BH�ћ�IE^�QPƛlX�T�P`��9%	U� ���]	��/�<&^�� �K8F�^ ϝ���oZ,�n�������B,�V����������l�szj�R�7��^������e�{�L��bd���:��S�#1��L��LB��Sƀ��1�l.x ���X+����ӵei](��+!+�X�I��>~/ww*\�L3Ş8Z>ǁ�gT��*ڒњ�>Q���wȲP��ڈ�Ɛű�c����|�YT�-�����)r����ʧ��9bs�xp��1�GY��	��ij@$�W��|�Pe��j}kA=����[Uic.U�#�lQH&���.ǎ��F��
������~�7��P\��o%��"45#[�>�$P�Z�>���P�>�<�����g���?�}�Ar��D8 }k���C�:���DӜ)e��@`P� "���EB3j%�.΂-��0�O�,��H��FB�82����#����H,=�9.�S(��7+R��=˙����g�Q���Խ�@��4����ޜ5��a�n�f�VU��a<����LE,�)
�t�J�0-����u�p`���6��]��Hi�;Y��⢚µ�@�l��)���]IJ��+'�W�����ld��W΂��w���5�9�<�_�SF�����e��:k��*~���&E��Fjgb��tҶ�I'�˖w2';l��5D�����_���=p�E(�����3������	���'�ۣ�V�3��p�-�z�qB����5jl��a��m�ET��ʄ�����=�iaj����?��J��Mb��<Ɛ@	�5E��I��b`ڍv�P�Wz�T��o��pR$�2u�����Qt�a
�ž1���w;�υ���y����/ث�@K1G�,k9�<}� ��<\S[���S^H�Ě�|>6`�n�3���V��|=�|����!8�ʝM�I$3>�Ԥ;ΒT�#z�j�ʜ�*�}�#�Vm�Β���au��N�_ R��s��$�[Y�i���Ħ��#�2L^�aDb����A�O�͡54nz*�����cN<�r|����:��xÔ����w�����@���}8�����~��匰�;�c�5W˖,�Z#Jcp��R�5��e�}h3��(���M�\ۅ��6������ �	0�`�A�0Z��\���VM����w=���l�o�[,ZhB��t��N���*�v�"9�Q��Q?�)�����^b-T2�P[���}�6}�����2�0� X�2TUGz�#q&ڼ}�a_��\pT��`��I�۲��O`M����D#q�/;��_�:�����+�7���d�%ul��B%VӍ�B}���PU���OV�����i$��ϫ?#���dtV}|M>�牒FG��:�P�3�T_���N�P*�k����`��ؽE��oeT�"��v:4nuW����R�L`x��N�4a�O^����͓�.\�	��L����{WoB�nM�_Z��޺�rcw,��F��n�~x�ט�B�W���5b�KՆ�t��L�\JފV�Z�Sj�'t�u�Թw�wZp�����=@�<ي٩
)c�u�J��}^�G31E��jKRR�y}���ݖd�d�l�ק����.���$�
�z�=�1fR�ȏV� @��Q���{
e��$�%@Zõj#��#��2����Mt�^)���������R.u�'�˾���PG��`�J�k��0��T�d)�,ڵ��Ͼ�-u��Ip�.9d�m0����w�Ǭ":c:'פ	3q(Α@�e��ѫ�/����緱7�h	��� �Vʵ�	�������D��-���T���䄯ш0�oz������/:��Z4S�+w��h�6)ۄr�My�}T�e����{�� � �E��c����&����3�J�>*Y\���������|��r�Į�S(�3�BA�DC�u�Y�S��˸�#�LF����ל�:ϥ�1�)h�B�Q?짢�c�Xq�����?|*��ZZK�:N�!�	�o��񠠻�r��M�?:����
`Zn�G�4�{���N9)o���C���e@%u��îPdK	��C{����b^��'�z��>�dZ�m��|^]{T�lΪ�wɷ�v��=k����������D0�6�w�X�!4�P���d�����=��	[��`Å2A�1�<�f���|�W:!��s��u����Z���V5jX�'�@ ��z��g`������@�����r��k�5��s,�b#h~��<�x�~H �r����u�h�����11�	\C>�qz�5�.���R�'��d�wۊZ��]ٱfo�^�I��^�b�3~�,�iO�룩L�_h���fn!	K�A*^d�ǻ�ǧ�xE<l�}��A�Á�f��7!�ь��<'�RoL���B8�6���86�H�鮦j
�B0� R*+������O$��n(�qh�CmW4N�3��{u�������X�əm�e��R��/f}u��2`d�;��!̓S5�1���6�	9�:v��s�?è�c��0��oW�`s�p�`�)&�8l93Ztx4�'� ��,���ٛ���'����ᙙ���� 粶3f��=�lc�<�:�z�=�"�Z��V�I�D�A$g��M"��Դ������2�G:���� "v��3��AE���H�=�L�"�(��'4��9�3�n�0҉,:�I-2����c�פ�dW��S,�e��ZF>F��֥Б
=z �ap<�?T҈��^�o:QGR����乷n����ͦS@~n�ao�&���5��mS<�i�A�h'w��Zgc����*�S�w�e��"�.h�|B��Q��5B��J�Eķ��}N.��݄�jn��8L��-uJ��6�fr�/?��y#�9�������=PsxIDM�ߍ%T���,�50��V��>έ6�鸷���ٚ�ݦ�b���ֿ^DusuM����E�{]��P}�>�YHYa��|i����Q�P��n	�P���j�\�/�x�F�Vn�	>�0Z����nmX��=�~�!�7,މG������ ,ʯ�r>�j�Q�'�����>���	p"��\&��N�MTX^���.�z[R�Fw�MJ�pV�˼}��u��+d�h3�(�@v�k���5
 ��� *�ߑ"Ө��O˶����6���|GK���_=]��p�A{I�����<��#p.���@5��d�"B6�zZ Pa���I)�R]�r*Í�.>���"����u��$�N�[�ĩ?�� !�j�&7���vz7̂��a3��+��?�$���E2F�h�4��P
�>U��<E��S'�kc-_�K�~G36wb^^LN!f��]r?�D��͂���I3����,��6�%����c�A��hA�� D�?��̧��1=��J����~C|�A��1�r��K�{uV!��嘽�����&Ҡ��}�����Xڠ_/w�`�Fg'5S�j�료�j����;s�M���I�a�wCDj�n9��0����8�����P�g���f����1X�#ٛ�B�p$����Sd�O���@�,��hƒ��"��Y��V\*`��#u��*P�0l�W�x�����.�fs�{�m�p�-@H�����R��7`)����2�w?�Q�oo,���g#-(��&�~Q>!�+16g*(�Nt/_qd�/����:E�����zi Nn�EZ�.d�e\�� _,�0���8)�PRk����9�]2�ؿU�� [��n���Q�0���)��e=��>�v���S�t�ϋ��)�,Y�ߋ�+t�����yCpS$�B�`�`
�uv/�S�#��q	��ٰ�Y�1���|2�r���vT�k��<�$���q�_��e?���E���c��j��Q�"1F��Ӕk���8�u��.� s�偊cf����rFC�D	5���1�A��t�L�'�I읯V���Qε���[��]�I/Q6�L�ƀ��|2K3�8<6Z�I=���f֏ɒ-{:�\�b%&���ΰܲ#
�O�kMz����3����QSh�^�v����.ڡ(�=�ah��@��&$K:��]�~%�F�c���)e9��ߺ�}7۪�5ac���`��zx���w� h����V�XR˙0	f������Q�W??4���с�����E�+x��Z��Y�C2J!ٳ�z�����E�\�*��@*��Q�դ�"ᖤ��*u�4@.E1f��l}/p
~���"_�V!*y�E�o�7Mo���v��5����5��k]�Fa-�@�q4�^�Y������}$�vei�󃑛��*X���T�o�X��nc�͞�欈������H�<��/"�[��9��,C��ʩ�1gv�n�;j��tEJ���6���ș<����dț���<S�v���E�z�td���VF��f��N�)��t�E�)����P?�9�R�-N޼d�	P~�7�w�גC;6Lܺ"bE�$�5G'�JB<�j�!�W�R�E5�K�8�q�A�H�<��z?ZSRkBg��)ȕX(i�+�-��}3Ӑ��M`�����m��O�5ʕ��ng�l3����m���w�������R��r��,|�K2�5���E�j����U�nàC �Lލs�=�OXVCss��4�ml`�3��K
;���B�M�tG�<�$�/�q��	�ͮ�v>H�Cb�CI5����=\W|\>b����s$��T�����<Ϙ� �#�o;!-ޓy���mjN1:&E����g�2SG���)�Fe_s�4�Z����~Y
��L��z�՜k��}Dj|P��߭�P�e�P@�fr���W`�=$��u(@�g��-=*��U1P*��6c�"*	� gê�j蔱nC!�­�W��z�ɘx~�¾�/#�����t����s�W��I�Dh)m�6	���(�:�����~Y��(���DQ�����zttY���l�ո���5�Zq!��Z�fp�x�v~ֆ�}X�e1��Q�ڿ=�	=	���W�4�n?�Ӧ��-��L:��"އ�2�������*~N��v��9��PQ�%ia���N�~F��mX���-��^E�UY�[� %Ke�����躐@x�+�[��v�=��$kv��¨�Ȩ�|.��6^�d��39�}D�Q���h�E�����*w�*J4p";��~~<��o){)J��`Uf�o�t���iӉp��׿7��LG"KE�O,E<ݡD�^�@����F����^�� Xll�y+��$����.�kVI�4����+�v1�6u=����S��p	B����Z� g�Sd�Eq������2{��
�δ�M2�|��y�$d^��*R]��逡{����J����s'��{���9�jr݁!i�G9���M�F2��� �wڀ���KZz��а}s�p�&�q����NI�#���m���r��ڦ�mF�Cx�.p���~ź���h�Cpb�X�@���s`GR�j���  s�
�9i;d�����c��qX���'e!��F�U
��n;�ơ���c95�nt>*c���r]��)FY���Uh��̉<k�#��T��)!�d��Ι'� HDLU�y5z��|łɂZht�D��Oj����pT��/8�T���*�c<lS(�L��w%?��Q���@�<���a�2�ݠ^��\)�k�$R�"�����2��{��L�G6*�;-��S��\P-�#%_�pu~��v� �p/���x��%�!�	�W��:�5V��b18y�����shj���OĻ�7w���j#kf���f�=��_ j1a��1�4�X���d��?*�3�$��D:/�NB��⩠����W^�3%*4���Y�!S�&H����y*�4�{G�M�ˢ�]r�}�,���xN��Î�l)�.�Ct�o�"ޡL��2	Ȱ�*���Q���m�^1��̆�+g��p��l���I 	Zql���D�_'�J��?�����%#%�p��+���I�F�01�s(%A�/`w��2s倇k��$��[�;CQ��!���
�mt����C#�QLc=�@��G��CЮ]�_P-��)ї, ����)KQ+P�5��A�e�rv;뒈��ć�zdƜ).j����i	5��W��꣝�x����<��b)��@#!~#�!}���Ó��\��!���8�����r�6ߡ��S�.�L���I@�VV:�'/�`�;��	����5@��alpyĩ���_����1�f@�(��3\��[M+�K	J�<�)*��d��&bn.�S�e[���+3�px�ʯ��8P.8N��d�0z/g)e7�IMJ+dE����z�?�]z���D�w��)7bɥ��J;Zt �f*�X���|D+U�C  }��S��ά�YJQ�����\Q��K���9�O�9`0�
�������f��ݰ�
�xy����%T�|G�և�U7���~�=x�@&)�h���W�n���lO�Ŕ��_ڄ���3ޔ�����Fn`�}t���%��{�~A��BCԍ5�!� +E�P�<��n�;��4N>�b��ԓ�\Z�T�Yj��*����+ ���E��
�%�S�e�	�SXRfB�_R�fx!��b��h�"NH��;��0t�S�('c�>�'ӑ��B��o���U�V�� w˧l������?t�b$����^/��E<�4��K;	F!I����6�r"�BY"F�麚e�f�|i3ixxpZ͘�4!�=��!���.��}��w^'�(!����׬X��x�y�|E�{<��f�@ڊb��6��=��M����G��[��X�=�bY������~O��0� �$�@�r��r\~�L;�"p�Z�?�;��z�]%��ic�f� �|�RM�/f���� ��j�XA]����h��io��w�C�� ����
+ϖ�hԴ��i��H~��%�&�u�~�ZZ?���-f�qCJ� )�Q�g�a'(nu`��ए<�F��\:\I�f��2];��E�s
.s�\��	�����oi6�T,p�v�Oe�4���Dx|46�%��dSx�|�m��wr��Ϝ<�ә�Y��?�P� ��Ϝ�~0E��S3���c_�d�ͅ�Q &���2�Dj��oA�������ШW����<+�<���-��9W�e��:h
"�W��\C?Wߔ��0���	�v�Q4 �S����;�@�~�wA59���&t��1�OO�0Lz:� ��9a� ���n�bn�
�N�~P�=�Ǟ�H:
7�ܦ�t��ˇ$�K�l��TC���j�HH�)�\�0 ��ҕ��F��Xa]N��x�G=MU9q�}�S�f�5�^��L$�Y�H3��>h�x�hd��*�m"!��R�*�`�ieM��	X���)��kbR���u�G�fm4��X�;1��b[��n ��j�m�������s�p�ӵ\�n	�
{�7��G� �9d��=h�l�$r�C����fkA�d��愅��D���ݍ'�Ҷ��l�`�S&�c�f\�}��{R_��{�Z�|o�#D��!����Ϋ������������գ����b�i����]��a�?Lۈ�=-[�r�G�e�.3T�\|�!9�)��l�1R{mp���x9t��9�K����2��[0 j����|V��[���� �ӽ���o4:[�:��v�Fw�|�����p�M�d&�7ڌPH�]=ո�Ȉ�Ny�V⼕�eW�`.�nN8>�ׅ��2CO=����\�:\��a��&����2m�B���J��J�Gj�1m�J�~�' +�*1�\q���8~��O�+�7-9[K�2����|�� ��c̊#�k���(dz2�2TJ�rk���z��`��3N`U� -j� -�3�(��-�=�РA�YZNT��[k�����$c�G�����9:mm��|�:���F>�����Z�)�1��S1EW$Tts�Y#���'���������hކoߍ��i�*�*��2�U�`�S�b��u���[�4�sرہ0z�aG��h�9R=Y%Zޯ����"R��!��{���m5�S����(j�p�rS�����Rx����#mԻ-S��	��K��������B^:�}���y3���ʻ�MSj+�"�2���SIsbK4���'�kt�AL���&��r�Ø�3T��9:��2��bf�6�G���V�0�Y!�{�6�]2��Ҥ
�Fc7W��&_�Ƈt$M]��ﺭ��gӀ��e8���@�������,��
���0�4���(H�zc�� �^��!]k�t��E������R�-���Y�Zz?6����+{wY"d �L���+y���%���h/c�CYKM�3�w��|�'��������q죊������ ��N�eL�%�g���M��ҍW��x+����Y�ٙ�7���9�7�q�?W��� y�ү��{Y��O$9�6	�^n�ŀ/hd�ֵ�ϕVZ�-.�:5�T�2P��[~R�`,1�Q�P�Hu]�?
�'��:u�#{��+y�T��?��S	ňͶ`?m8�@t���~-���hK�V�Uv���^�0�/^}�Yg"Cgd������^:�ަ&6��;�Ua'�Y¡͘�*~�#�cҦ���>���3��_5�繬�ZXy.Fɵ9�����k�g��s���ʹ1�u&U��ho��-����g�=�?�Z�����W(��l$��q^�Y#WQ���Vߞ�^Z�+���\K�pC�G�Z ���Mn���?���v$������9Y5���{s���ۋ�r���t�1�rG�����5+f�3NBw!�D ���{��ҠM�H��;S�(�Ž�����"\q"M�o+Љ��n .�:c���i�I^�3��&���=���{�9��o��]��ǥ)Z;b�C�W.���1?J��O���V���9~$�����+�)8L�B�)4��0�4�T#Ќ����ZƵ�Ba=�m�# ��xd����9hy���$9^����
� ��wH!�&�^Π ��t,5Iߴ��4[�bp�C����ȇ�6��&Iy�%z�X��O��1%�#�$ˠ�&��P�J��	_'�l9�$�d3�&���,W�O�5j݀��-�xBI�^q_�,�]YmR��a� ?�J��O��8���"H��Z��ͷ��ER`A��3�El�q�����7��puV���,�Cx��n, /���`���^�fE�Z�846���]g0���虞�x�H3�՟/$���������To]�h�?��Rz�p;`΂_w� �LUϻ����P�����c�� �X��Ywn�؆��p�Zw����|е`�-t��	;��p9 ^p�~���=x��K�^��(�fNb��6�M�B��lh��(��:)�8uI��A��*ͧ���L+r}��ߖ0-�y�Q�nda��̎q�/���1|܈}��׳R�ʱ��3[�˫��_:��n�{�Qk�Uc��'�����͎7�>E�:�0����@0J���7�v;���0&��vJv\���[ɤ�w��|�wc�I�Q�Sӯam�T1��l�$
x��n�����a<���;P���8������V�|��w"�
��ٕ�R-G(N�;
�N�^��q��4�,��4�t���@�{H�K��ǥ���.���>�٩�y���;��8�H_BBI��a��I�y/�t��]��v@�t(]̯��a��{
?U�l!�*X�(��W��T�,~6��X�}.�I�>[C֌g*�SUyDH;�
݀�^6�?,��+�w1�,�uh��,]:���f����_��g�s��q?��[G�;�n3��L�w���E�xԼ�n�=#�#H��RQ�d�i�_� vi�jp�����s��8tN"�)����T�	�F�>óe�l*�_9�9�����.|��~i�ý�z�8"E�̌��d&r��1p(k�8+�}ƕ��p�;���Ik��(�':˂u+{��;�,:
'�7�`�*7=��p�C��$��1�J�S��y�3�a���a�@0:�(H�q��$��	{�<"��Ho�Ky&�D��*8�~ͺ��	�����ؓ\�e�������({����i-�(��m*z8�*Cb��K+�e  7�?r]IR4�Pm��Θ��ss}���S������v�,8�1q�ܛ�� �>9�K_Տ�g^���J��A����[��I���|��Y�Z��JJ�|�΁̝��S:޵����R-��h���%,
r�(焉��s&ꂵK�`+^Y!���\��o2��&`\�:�i��fb���j��eL�k�N*����3}ץE��N�UӚk��O�Q��?yY %歕cv��H�wj�@�bunօ#U��\�ύ�f��?k��(�:�IU�R����V�ܟ��j�I}z�2_�g`�����J�ε֕�B��"�T􎐳����HQ���� ;C�<Z:���#F�mI,j��()1�J�@X����������|�=��1���-��TKp*�>��r�_��uxc���4�¾Z=9wtZ����G7y������<����&�L'��3�<�z
��q�i���y�<\��W�Z��_�S�u�n�|v���;n5��[3�`�}��c���͊��m����u��2ecD8��ǒ�����B����/>��!ӯf	�u��:��K�u�xU�!����A5Q�N.k��~F,����<��E�DTsSP,����ZWco���2G�l���X�l�j�*��O����P�S�#�����q`��5��͂��x�ѽ�G�E�
җ�s=)����_�\{��
l���ӡP�Ƴufl�E{ŝ\��Ӈ8m���˭�����!+;23�
����:H�$ҽf�f��g�վb����A<����;��p�+e����|v9�j���p�b*���:��[<��	]eZ�/��H��})�	��ㅣ\h/��T�ɜmd�O2��Bq�D��5����B6Jw~�GK�g���I��V��� ���C`8v�#�r9��V���ޫ?M�.x�����{a��@���Y�}���R�+ ��9����R�<��ov�؆nt�M����;d%?�<]kԢ�obMW%�)Z��<G�_�����Ӣ��
�Ľ@T~�<@�Jx]�g4�qs�.7whS��(��R�<�a4QZ�x���YW�
�e�*�817��h������cKQhDym	+/��: ^�G��S]�'�"P��~kD����3ћ�>������b~�3��j���6�RYKR�hf�{v|��\���s�b���	���#i��~�ş\��e�����m&\��'���}a���o�M��gxCkt�g����`��OW�ǗD��w�/9�–i������[�g�R�����Q`v���1�Xiʅ�t�Vd^��7�`{��!�O7�>W��ͼ!�i�m��S�d:���|�f�z=��G4�u�ÛG�����S�ډ6��qnh9� go[��j{���*��/�|���]�ܲ�����h���c��_i�Β�T�K"�c��{�2�"�:��&�7��̱cam�׭�jvBW�T��O�y	eJ�\VF��$�M(�5��7Xd&Vғ�/��SG�c�%M�U��N睵D]T��w���I�!$B[��_�`��`�ר�?X�9�4��a�ڈ�l\� Ji����;����6�![�26��>j�!%���m�X��;d�3(��}�#������wm�S"�0䁚��L���ħ�ܼ�G ��3;��E��B������y�^BP�Eg~��ۚ�iy�n���ɚV�STL_��($-;|��Ak��<�_���W��Xz~s��R��xeU�
'Gf����Z�wȯWr�6�??[��{�_��b�؛���P��̙��9HC[�O�&ǂ�g�{H��p�U7�[�~���n�h��Ɓ>�m����:PD�NY���q�@/��E?4t�9a�;/s{�Ȕ�7��Vޮ|z��?o\	_��pn.G`��#�7Z�'�r���ŁL�+�㻏��ď"�����]�A��MJ8[�k�F��,nYm�	$��B#�8�Fm���j����%:�Q�x뿻��M�f_�y��n��
���V���x���k� v��ȃ��i��Sgu�]m��xM��+����wO��O^�`�$�����h+mjmk }>/�`h D7����I�w����0/��k:J}��8!�- H��va��������i��eģ{N��Ol��+�+�Cl��)7<�:m����@W�O��/���|��]����^mJ�/���a���[�L���N(o�K����3�P��&�~��):���C���ݏP#TjA�luk�D̲+1h����,�^�Ԥ9Űu�ܒ�2��*��&���7� � Uw\������'�,��dg����$�W�.ľ2�>� 2��#�4S���C��mh|��_��03s�Q�iJ2i�o�"��Fc
:2p��z�F,슕h�/��M*��ԅ`�g,h�?���qU[D�%4t+ ������a�u��G��Z��è�ה�nx������Vy�h(%ÿ�1��}��6Ֆ�p�'��E�UU�QE���ZEP���/�,E��'๞��i�U nf���r�iж.q��x�4̌�y){�P��;t��:?ܤe�D��r��ӟ�ǻ2py�ÎKԻ�����c��}_��Ď��X���0�n����q�X��A>j9l�+:��	52��Kd�h��"tg$�����
Rq�.�r����j����%�&�dq�a:$"�j@O������%�v����s���*�Y�gL8���&[���R���2�`)�h�u�-線?i��͇�%W��6��l��{��)Ɖ;���[�~I�����	I )v����y��6s����=�<	� ���-�f70@k�g�N/�JY����$@���u�x������d:���k,�H��Ft��������>C��k��%��|@�o���m�d)���3�}Lϭ??�����%W�FՅP�����fVӚ�n�ohE��R^[�IwD�t��)%9��B}x�p�emi������k��+7�]OshB�)��7������?]���{Eƈb�M�R��P�����+��n�E�9#Y���Ĥ�|�q��D2�m�BH*.�� Y�B� 8n�HO�;�@>�Nĸc��r`3���;�\#F�v�0�����C�W�qh���0��8���N��E "=X�t
�Nz*֞@.4����:+�P����ĥJ��o�yw*&�!y�*ƶ�J���BTQ���g~>�D�T����D�ϼx�/��\e�e_{Qt$D"9��rZҕgvz�1���B
�#im!ՙu�88��{�L�/�q� Y�����Yy����'�@n�m���I�^IR�&e�onkP�u���r;���:�qqf����Y��6�%wj���Hx�@O��cR�
#��(��ǖ׊�a�YK�:�P>8��,'���p�K?��ߵ��9�$Ld�B�cz�g4�v��(Ċeg�����I,�ͅ*��[����a�MFȣ�zY �.�~]@s�٪�QL�m�V�T:�1"���80�n�L�ɏ'��Á-Z�b_h��j�(UG�N��v�a��r��*��1�a��*�`+M����!�$�D�諞{ G?�=ȭ�t��20���R�s`�!q�NXMc�G�<�|�; �� �]�غ�V�cB=^��h�8�z}��~]�c²�K�}�/� ��zh��y��0�����ҝ@PAMt�Ï[ڮT���̦q�a҅��Z��*��j%g�-����y7��w�g��X�0}�.���[uN˯�ɑဎ���|
} 0��ވ�[���;��#�ζ��l_Mu㞻���ɀn� ��)4��nr/T ����+�bz�V`?�������(;���_L��������j��|%c#�m�*N^��.
�#LP��skL��"���p��{���%�������]H�D����b��Y`3�O}�J� ʅ�;�X�}rQO�]o�'G޾��Eb-�*���� �Y�Z������$�����CC��J$[lUf/��0Wm!Y�Z���<���)���d��)�Y�G���������P�!��/~����7����c���TCop�����{i��L5}0M���N'2�	�SFMM�e����� ���N����h�'S�	���E�<�f�N>�4줝,����}����>:�%�a�y�źԖg��ԃ��/�ʙܿ��[�03�Չ��2}xk��󠚶AЄ"a����T�*:��/>���8K�ɉ�K&�p�*#I�Zc��\P~���H/r����/�g˗����.�DM��)W��w�w1���/ ��|+C���;����}$���{�'q�r��8��P#� xN����hN�G^$��|��y>��N�lu���:�������y�&&�G��Bh{[d�z^:\���F�G`�/w��� �B�VEe������b�V��(��U�k�9ڵ$�r��sI{6���E�\կ�n�oSl���,�� 9�5�!�ƚ$��FI����4�G��۟xQ�nx��X�V@A��"��4��G�ѹ�Ao�6w�Kc|pp�y+^�[i���)���R�ݖ�A���Y���
�͑�U��3�D�xI/�F57pdߙ	���$��V�S2t����؏�h���Y�f���L�0�J��1^[� Q>���N��r�d�Qa>Ҩ�E٪$��k���ǍH�7��C�dq��������E��OPk�K��%+Ŗ}�{�S EGUB���.z��CQ��[�F����$��D��'4��-���_�Xњi<��� �B��Ć�;nM&G�)�یc-4��V͜IpS9k�`��"+�*��!�Y��Sa�K=�j, -�#qܽ�_&�Lؗ��j'�D2�
� ��-\THIN�ͪ�$�"�"�9? R>G�<��������s��.xt1�`V�c���~��fN��0q�������I��lpX��Y�j�#�����ۣ��ȫ�Myd���+�pO7B9@�]��lo�eV��l�B��H<ҽk��q�^?����p���=�D .y����
4Q0�_܌�i;ك$��e	w�2c�/���u���hT�!Z��{�dJ��u���51�1]cCh�Ç�t��4�Ŗ�hđ����}S��p#�G���cMObۼ���� ��P�%�A��N�m�����xGp?����׫u�ҧ3�ؒ�0�t�B���J2O�o�}�z����J�;��q�����|��q��((�c[��@��4�X�9m�f����V��	�*vת��
��jX�*c��jE4떀�<7ʩ�Q�*#*zJúpCFe�Λ��jW׆��v�+檊ʊ[z�)_����%vS�P<�Bzſnx1qh��Oq�c��C���*�%�P����d�ږ�Rx����lP��%�����mIM��M$�R�Ƹ���v�?�ءW��-��Peϗ�'����-����:��ܮ�������s�	'%覒]�5|��kR�Z�i�����i���ؑE?(<��m*[�,b��F��Fw�)sfiu��'�g�����+'�$'�<��	�H��� ���"��v�$[�(/aU)�뻰r =��6�f�_��VU�y�a��?��^2��'�mZ�}]A��ɳ˹�6(���5C��l�Ӝ�m:D������$�F!yM/c�4U�C�q�A��=x'�y�5��Xs]��ᒑ1خ�t����e�(�&�L�x��=�p���3k3��!P����t>��'�Vo�w�ڳJ�z p��C����������K��4K��#%�E)J���x��G:�t�=��X����FE��]~\���5�9\ܲV9��INT3Q����:#b��~�~�B����t��
|8e��m�.�0�Ac�|	;�jU�%~��C\�3)��^f�/t��t<iD�H!-v���ʧ����L�=m0������	J:Aϱ�Df!���פS̀��3��:ۦ��u���x�VA �ܘYך�a;W�K�`N�:�d9�ð�}x��3�^Q�Q ���������q��6E���g,T�6��]/;0E�����u4p"��&��>N8��N�#Ќ���W�Z[�I���m"�Zc��}&5pTWP���ea�g�
=�:�0$s�I=#JZ�D���Q��
�z �,�;H}�_�$֧�/��7_�w c$��!�
�����&7�P2��#�6��ʠ1ݼT����2�f��v��OU)Z�����Nn��k�i�±��ZÒZb�R[��M���8�&�Ʀ�Y0��բnh�U��/�����`�g��*ؘE�o�F�Nݏ��r��=Z�����p���4���~��v�Z2CyM�U�W�:�'J�V��U�1p� 0ӷ�͂~U<��M�ޯ*/��X���|�S�W���������IE"J�12�K�d6��h@��2�����W/����T�*��s�1��ɮ�\p�Y��ľ�= �LaU����}�,�HS�	HPi2�Z�	t�	������-O~���Z?eGh�X�Eg&�3Gv�ʸ�����õ�� �d�3�����T.�K�CU�:>�2-k��w����?1�02W�T��50C����v�d�E*��ɵ���̘ADH��7Dyq�4D˟R�G� ��9ģW���i�D�m�n�X%�4�����`I�դ��h(7%i{�HF�d �y��ꁩ����h0Bߊ���h�,�����rt�]�%����QU�@�|�o��ޕ��G�~��b�kN�*��I���S'@�`R�	ǥ��qB�E����?�xӷ�;�3��D�shQ�3�CP�G'�<J�O��9Z����~2�'�$H���C=x�䨧O�\�h��+��Ż�T��r`��H�f�"&b�&f6�$ ��aJ��닍���UQ��Y�Lj��� 6��$�Qq��(�M�����P��c���EX�Zt����B�U�1-P8nEK*��@E6��m*�uч.ЭM7'�o5��!f/a('�Ą��T#,dܹ���$��(����f�.�L�DP�r��r� ��\/�X�eT�=(7X�4���7%�������[��-�Y�9�S^����.1s�8>�L��X�F�A�y��SS�d��Y�g�(Ъ�nd����Ш,���	�"}c@Z�_���w��5�#�U6$�.�ٸR�z��7q<�>��
��9�6�C�.�H��Ȩ�,�����N<"�*8G_=�r�H+����7|�>���v�2˰��U�Qj������0��`e�����+fe.H:t���sGH|$��K�r�wX}�d��#({#\N�1} �_O|M���\ �y�����3�W�;e�8z���?P��np떊�.l�P����u�/-j#h�M}�7�`����,W}��V���p��l�k����~/CRc����'2�N�W#jq�~�`������m���y�Et�~��t�D�Qb<��Xi�.6�z8�5�0P�L�el�ޜ^ݟɤ�Q�j�%�hWs��$5#9�T��H�?��C�da��w0��!��]쳾��Y;�1_믷G�H�ĳj�ARa���QǞ-}��S�X�쀋�U�$^'�-���*C������cE;C=�f
�%s�F ;r����&�np4 w����ފ��1�B�~�뺾��8J/���P�ٺ��Rk¿�x?Q4O-W`����=g%�}��dS��u�ǋYI���X�x���|�c���`7�)��[DfUB�J�R�0w�0��&���g�Z϶��gt7!#�έ�Hݕ�1<�I�\�3��_;��xa���m������E${��󽣅��)`>r��N���8�J6�8m�CD$O-�;��|JUX���Zzќ/�8d��<�m�uA�	RX���ֲ���&ok�N��(b��Kt���+W����;��$n+x�|��i�9������,�^��ռ���~��c��4������k�d�2��[�/i�f6M��+,-TB���;f"���3�k��"Z'�,�/iI�*�6�z�A�qմ���f�z���h�aH?x�t
|B�p]Zjj��� ff�(�����葾��]�Qf�Ϙk璉O 6��0g-�9��&�J^��+�3�%��K��xvY���&2�Yi�Fѫ0��\8[\��,�c	��>hi�Z|/FBN!1���GW�<�Ǫ�ٕ����N? �6�6[^L��9�\}bd|�V�ǰ���t��>����������.�B��}7����)�O�N?����_I�y�L�
C��Љ��D$���@S��w{b	sBI�G��܁HZQ�������\
���9�Jʞ�c�~K�N�q���FG�$�b6`�Fw����X��.���B �6��9	���=N-3:���YAm�+�W�9�0L>�n$J�Ds��2��k�g�5K��] &�M��L�ک�(�. }F��a-M�#�^w%Tr�s���7��A,Mk�D9��~-F�����������24Oɦ��:�);������թ�2JNt2��wO�h������B�<˕u�����?�9���>�z�!���w�Vi�d&�8d�+MN"$o_h	�R7o�<�v�L�+���-����S-�ۙa��t|u�J:a������+LҖOg� K	�-����?�8Ft;^=s��45�*	e��
��VX���DV���v��in�C�Xf�L�Vؚ��ߊ9�E�/3澏�^on�a�8�z�U��tE���V74���25ek.0v�v�'�_/����3X�Q�dq;���8�^�:���X�mˡ6�!1|hC[k��lmK�!�E�>��un��A
��-��	I�69�*�ɼ�&\e��L����\�E��?����2U<����qr:�[bکVi!��P,(��-:߰u�}+2�H]\��%�O��̫C��<�MƁI�Z�jD�0��\Ioٖ��=��f =��f6<_�m�qŔ[j�FZ���3Pz�e?������E'�=�^?��vO�(�Q���=[�A�ohl~<��-�D߁��$w!&S��%��Pò�~��jj��K�DU��eA1+�	�`2���{Y@��O����ެ�������;Y�ynk$�b\C����o'�� b=1�Q�)����G���K`fi��C�$��Q���-1�'c+��w)�6� >mj�ٟy($��(���1�2|���U�"�Ą�
lL��;U���J~�2REU�������-�=>��� @KF	��as�y�j��b����
"�u�]MÐi���I|H,+'TԳb7{��'� m�;S�ik]��5���=����/��5p��&'����7�HYX��[>µ[��� �l�f�Z��֯���VIdG�2)��(�	[c���~�憐,�6�z?17���6�}BC��ƑC��;�I�},�w��G.��]xnUnGp{�oG�׵U���'��X��#� �M�vO뱛]6��^h�x�W� �|�M"1Y��i�b�;~�!��&�{�Cl��A��{$�s��=]=��+�L����Th����3"�\[%9���C��K?.wP�K���D�����6��R���[���>�b	~@H(��G��`4��iD��d��t�AcK���7�P��>��r@|5��8	���)ܴF_u6�� �?�~Ch��՞�Ռj��VR����AH�|�t'���tRΥ���I_jB\�]D��5sc�~Jm��"t�;�S}t+��U<����9��e���v��T�u�K��d����3��?ª v}��z�wT���b�L�7�\��ڳ6pa[~bܛ~BVCŰ��!��LN6���U��A��4�Wm+� �/�K�����y�"��I5
�� �s.��/A�\'Av1v�*�J��������2kl�3s�
�ߠ�T�Ň|o32Zl��&�V1Ϻ��0�!�*���T�a�ɀ��OA��Kֺ�0|MC�.����g���)�~������z�	J�&����u_�LmKxJ5n�'C�A��}��Kj�h��~Tг��/�1E\x�&�H����w�ݎ]&���k�/����{���V0��x1	c��Ϛ}O�7������&�fk���Ҹ"ə�]���p,��j?�ArU#"����`��J�ȶ�Z��f񱍜�<�YB�vA1d��8;�ue��OL�ɉ����%���i�}����H?S��n��ӑ�/���7���A�!��I;y7>b��ҩ��ץ�a�Xt�@�5T��?[ڻ���\-P$DF�{��P=S;��L�7敢2��W;CA�/��j��s�ԖO����?r�����_��`�.�ey狍�{϶G
0�����"������zi���=����(��Wۿ�#B������z�mI��2�83�Ϣ��NE�#:��xV����3\�q��(�r=���P�ͫ[���aaD	O���S,Z]f�{1;��IÐ����ɉ���3���4ܜ�s��[���p���M��7F���ߍ�r\Q�z���,f�2FRWxx�nȢ{�~�oB��FmO�u�S&!j?���*C��: K���Y�V����
#Lf�k��j���t���h�h$�AV��&:��8?&@I�b�8�bM��0�)5��T���D���MmU��vl8��w{���2�8������A�Np�-4RB�U��}�iM�x�.pҘ�["!:��!/Q�݂��e4Z���}+��cSď������A�ִufA��	���ɈK�v�[�k>Pe�.��Bf#�ȕ�t�+|��J�Jl_Y�3�$�/��
lg��:��+�C����,�b��~��I0 n��e�
�TS��ф��wZ %cB�Oʙ
�� w|û}6|���M
��8,�vq�����A��AL�
t��1ra��KX��y��o���6}N���� C�2�v#�4h���ؼ$���s���1�$Z��8�Q�AR�@Zi	�nB>��%a'�� x'��D't��<�$��f��/J�H>/j�)���'Woe�3�KS�F�����+Vѫ�n����''=v��>�����$�Y=���b���-VX�Zэ�l�sѪD��"�DP#�j^A�<�������� Zዐ�F��*V$��wv>�,�L-ah�����a����v�TjsU���Vl�7��ڤS�F��:��`������-�_Q���+��ژ�g҇��*1��T�ɉ�/L�-��[­�S�ulv�vR��M
޾��!�
uD��D%5T�A��0n8�o���>(Ϩ8��'�vŅ8`iW���[%��bĒ"���=!_"B���=
[��$ ��Ss����h\�
5,�]��Q�1<��ʸ���|KZA�:%
4�U8lZU]�x���B3�g����ߐ��;��ULib]9�|���O<�%�eQ�=��Ɵ��Q�	=�*��5��t9L�|���<���<�=tI��1��������h����0�����8|B��Y��[*�h��2�Ґ�.����>�1s�6��΀GɁ�_��eSj�[+��ǃ�����k��~F�����kO�M���ڡuW�0QN7s�#9[A!�@upU��4i��x�J9 ���^ ��g0�5"K
W�T�Bm�;A�9���.��յ�qƞ��[����ʿ���Dn��h#���'��A��ޯbȊ�YסvKop�:U'y�C���}����I3�-"
����lf��'a�0wl��8�q}2���]�,Tc$jW}Wj	b���ʱ��;|1����2e���V�7�]0��@��_���C��OZT��osSA���:���a򈹥��6��XG
-)g��~�.l���!�	�@:�
�B��h?]�/\�P=�ޫ�0�J�2,x U|8��xY��rj����,�X�O��@�:�c=����9`��P	;T$@V�o�]���$���������U���(���*�p%�z����9��5�b㳗wr�U]�t7z�3��&��\4Q�Ŕ>�:�%,-���[�3�����O����>vO5��J}[��ڴy6�$�~�#�Pd��Q$x�U>��3�l�#���M��{�^�Z���G�a����΄��3�No&���8<�q�?��m��0`��bh�x ��q%�鼼	��Uϑ�[�ߌ�J�Q��lpD��l��������� ����6"F�b�_�I��4>�=�3�����Ǒ3`���߂�ԋ�+V'+�sE���"/{}ЉDe�b��r3�)�S ����Z�&��Q_@9���o���WYY(�8���V8g_�rr=GA��|ut���?�����|�y'�qܛA`S_-нT�-62���?8�Dg̎��X3��
˦t����߶eֺp��]]:���H�h��p�Sy&zo�8*6�c �.:Ep]it5�z���J���9
���(�CΦ���v���o+�%d��6BtIf�t����f|���R��o;�����m�Z,�j�|�p�;��hZh�*��<�o���ws���MA��X���E�4��� �V�!5��bܶdv���R]T؜���e�^xO�Z���sIuJ�Mx�ؚg�?���U�ү�z�.
�v?/Y���1��=�R��;Erծ�=B;�w���]���K������Q����H�Y2H2x��4ӥq{Jx�][��+����`͜!$0������cs��xK�ʷ�_2kU�J�O>:IF+����7��ZQ$��+����ۤ����,��L:A�"�`��a���.��i�=�t`����g�.�}n�L�mʏ�.��5&܏��dV��6���ƍ���J0�_��c�d����7�����C|P_�>���FC$#�j�5�V2��q�er[~ky,�˜�����K�(qM}�^ysv�<l��E�U��->�q�%��&i�h�И���z�Wt�u_� �e��q������( ���c@�A�5^���\CE0��Y���� [��=v�W}y���S!>v,_"��G������s����2��mU)wm�!f�/I�E�)0���!
.�I�����j��J �F6(�.�'�>�V�ZUC-9�CZ0��e�:m���qZ[���0a���zH�A���O�A#�+o�#�3aT;i�R9c�o�)x�:˜�����[�C{��ɨ��hJ����2S�2`�=ِ�W)��E*[�Kg�	pv�%u���� 9s(��V��~�hNg�H�=��׹�_'���,�k i�,�Y�_;��|Y�3�U�y��/���f��h/�Kd����s���D$�r;~�~�v��J�߫vض�;P�r�>�I�q4��#���aO�;4�Vms,տ�)����@�M�3��)>Y�-R���@b��Or:�}�	Q`����? }q�w�EK�E���%��-�n��Σ	+]?X6@�J,��A]���
�ȿ������}O��om^��E���?���F�����'�5�B�m�K���9?� h-�5�%"#��I����Z��g����蕅����Z�=�!AX~V�_ft�^�i8\`��m�T����D�{5���t_ќ��}�bu��C[����ܸd߀��r����z~r�51�A	!]2�\=�N��j�8���f���9ϼ.���h�е�(�h�~�㓼|:^���d�j jKl��]B��՘���g2�M��l��Jw�*v��/��k� ~�w���u���y:��/d��f��TR��5 q�(�B�3���ך'���#�\�Q]U�Ɠ�@3�Nq$��Kz����~+�t�`9�C�۩\#��~���rY4N���d�3I����ѐ�t�=Zy��(�B'�v�������tY��>pP�!������у�%]v�� ���a�p6���^r�M�,�1N�X]��f���� ��G�JÕͷ\��EGABg���u|X�J�m.P��1ql�o��t���G�Ô=����b^��'&I��7�sp	*ξ�
| ��F��W�)]�Vq�AQ#[iAU�t��g�;����� +6�hf��N����z�p��.�En)�GXx,���̉��f9��4�5}�ܯYB���<#�t��c�cms�����t��o�(TC5��Nd��R 0�(��
Z�����F�ڋx��v�⢯R�=iX�|)�i�G�Uw�<B��V	�
�8v� `a7��e6����MK�X;��t������յ��.�H��<ɢ����.8K�Ӵ~R��q:Mfu̿�j����-u�$�ib_]��y��� (���s�\�
(��]T�=�ý��e�'��[U�C��g���l�`&*��5Z��_(�3E<�}�0(,*��~��>�/�g*�b!�l�Xe��/<�����x� �S���ʌ�<�h� ��e:�?݃�O\�����$�]�7�eцo%��kꭁ!G%p����{UcIӷ@9������/���IȞ�����`�|��J��,�CtA�ik��W j����5{-���|�Z��y�lޱ�ɋ���#v��Ff��G\ѐ�I^(�@K8p�Z��rjӫ�$h{��7)#�g2r�4��5y�T�Q��MT�M�ʆ��w�PL�qύyT�eI|b�T��y�as�_xV��0���`�`w|4*/���Y��xz�����k����ryO
m��yNyg�?1:~?f]�9\On.�7]�	�����a̼V�����ɑ��wG��-'�u(3]Y.������+H@�׾%�0S�VQ��ͭ�t���O���/q�������L���25����-��@Z�Ի�h�E��:�rƓYw!��C0��IQW�.)�;���$�k,#@@"S�(��arE �RڔNb�� wC;�ڽw�_��PMލZ������'+,���N�:�JR/i{5�6��#�D��1m_�rk���R�#�<ZNҧ�2"�e���>�m��*]�.ȃ|�����9�p��5��l�������>8}��v8����ѭ�?fa]�[���"��b0���Oyc�Z�t+W���fC_<��:� :�Ŝ�����Ľ����Q�F'�茷C8ܱ�ָз���(7�IM����8�~�(������v R�¾�d�xkZ�Q��lGW����X���VI�S��0����|�E�d F3]�;�cV�[ë́-���ŝx���(�N6^��u?~�s��+���v���T��3�f�U�UN�W�!]<���L���;��r�O�u_�����G8g�@��r3�@��R|vo��_s�>���R(��},.�j�Ƨ~���/�/YF��+`�W*P�^
��)��lJ����t���_je�u�;���bϝ�,�6e5!ؚ̾��)��bMOC8���]|��1��;�D� �����h��}φ�|?X�L�y1��L�u��Pa�K�o�G��zsJ��Fv�Ӵ��KȂ�r�k!��G'�d+ cQ�D$����H+�m��f�n�{Ѥ�Z �^����Bm! �۵t&��qk��M�7�In�|CKk��~�8�H�PB��=Z��E�
�/W�e�BKǘ+��i5��\=���=������+!5h��~� ���@ƍ&b���hO��k�������ΐ�q��;L?(�AZ��3�nپ*���{���m`o����e O�)U����_`�����]�W�=��Z�
+����?L��zΰu����=�u�vp�A�<�F��q��Z�E��8�3���YE�����/���(n�U�wܚ�  l�&@�WV�I���S���H�V��*&����>�=���k� !&�:�k�G�E���>UP�zĭ�a\�=�=22�x����)����̊���-��\�x�����>��"i��
R|�;�0��\�f^3P��raX��V�4Ib�AYLU�?h��R�ՕD(��P
&l�q��B�&]����O*�.�F�B'��r�٥:���Zf�_�jo$�V'\��<s sAv ��ɢ-�5e����b�Э��75�3s�m�����O��J���0?q�N����u5%U>�S�/�[��K�/�~�u�N��'�U�N�<��h�J�w��E	-�_}m|t��2��ڟ.Ց���`e�_"Ȇ8xz�a!͗Ǣ��U�Q�<I��`��v��y�l՝}�	�n�>���6�+:��@Wc"���믏ّAg�-���n5��Z�?�r=ᬍY� ����ڜ<��8��������M~Y�6MQCKr�Wܯ+@�6	��>Hth}��1&B	v��oh�uH���ǣo�>���	��A+�!|�zNˣy!m���7Èk#��Q�*~�g�v�Zd~�E����~���Ҙ�i�*�����옍�sU�N��+P��!U/'��bT�5q�:jmB�(�I�G.���	��M+]�o�j}Vm��)vKkl�5�`±�-������R�@Yb�����Cub��%�r�����(�)�\�\]� ;8�������%�4@>0,�}���>��A5O��f�
Ǎ_G3֔��q뗾# �
m����FR�$�c�x�܏҇i25��i��I�l�T/�'_/>#pN�ja_@�e,D� ��ۮ:��џ���m��L���
��>�x
��EY�����?mR��X\�ݖɸ6�}2�W�g	E�~s�m�e~U٢�h@�Y���0l֍�0f�(���bhDP��p��uؙ#��^=���vDo�tmc�k~���J���D�3Ji��w��BK��9'��g}8�l�a���W��\���>@��	��,Q��Ram��e����B[.�\N!o�/�J}{�^�<����˂���eZ33���M�=h������n@#e�d:��G�T�~��|7Zv�׷�HFr}� c؇O�;� �n##����(�&.�kS^��LqB����TOM4v�c�R�1d�&�uH!ob��'K�0H�V	Y;�ٙl�d޻$|��k\��i�<���欁�O���(U�(�>��[X���U�� ܇¿�ʁ��(�\��������Ӻ�pNi�>O�mSh'��71Ɨ}#�"!	U���Lbn�O�� ��.���x���Y�������J��H;i
�!z7Pԃ�1.�ɲ����y<� ��ZŻS�邰�ª�Ŗ>���U���;��J�ի�m��kD��G���]F̘c`
q�z��X�a�w��?;��G�v,���
�L!p�����Yx���Ir�Drep��e�����k�	[]�uN*_�P����Z����"���>��\�C��.�.���3Y���O�9-R�/7��ٴш���%{�(���H��hw��	vk�T��Ɂ�$�:_c(�N���\����-��3l,6JTp��V�ۋ����;�%�?m.7�Ҿud��@�x���W������0�vD�L������2��e�U��q>_�R�ВO��Y�.؁tB;z+Gi����}��@�s��e�>��d.^�E짘{���s���t���m�Y(��A��c�a�z=w'8��^%Mڏ� A/cz%�n�T�D����t�K����q�����ά����'�7l]�p�cT��Zj��J=���#���8��W��K�����W�p%�zV�<���U�K�Y�2g�:��3arF�@3}@꘏c��rƆl�ΘwF�"�+���=�)ꑩ��,'8��r��2z;�c�9�}n[ԭA�k�M=>HP����`[��t7�#')��i��&r�I������%��(�4��F?c��
��O*9�	�E��H��粷�⣽~ m:T/g9{�E�Q:OfSur6,J�q�j��ե!׆[ ��ENVFJ�zD.]"�ʧ�D{���c�Yŵ�̕_D��>.i?�͢|hf���4�U5prj5�������RE��ۆ<C�u�FuF�d�C5��5Ɍ�[�'�<^�w�[���o�t��UN� j�:���9]\m �eϚ�j���H�r��j��JmFؑYQ}P&������I.t_��t��j�F��8HTB�!2��&��W&xY ��KF-�YO?`3ar��]��SA�u{��!J�v �$;#�Ѩo�cU�=
�W3�u:�?^�xG��q�C��	�j~q���<n�6��
��@����Mc�ǉV����l��a<Jl3����O���$Po�`��"~���`�'������N�&g��t|\��P��Jj�^��$.���_~J�����B���)���<p�Z	]���E�qQ��З�Q6v�x>	6?��垩�?j7b����v�/�s����[c~^܄�9��Lj��ȍ�w~-����7v�6]�B9i�9+��- 6�Aj���u���J�\��Ѓ;�[}G��|&���˼w8ba.ݰ���{��������Rű��f�����f��Cv�i���B��L
���Q%�;��������V�@%�5��ڀ�N:�i�%�Ī�yM��9PtC�hp<��_��x�xK�S�着Ft�+'����b����M���|�����ӻD� ������Z|ɚ2Tk�e/���o�'��=���T�p�D	EZ@iy[�RS�|�T� ��m�pI,j>HD��C4��y��T�\E���	�B�<�
4UsKP[.�U��I�T2!�a�PTZ�u��3�[��(�Q^�=W?Ge�8�e۾;�5h<��1��!K3]	н�ǡF�,*����n��ED���5m�_*e�.U�1�X,��r&��.zO���x������-MQ�e��_K�E��O˧�:�[�i�e���tJU�>�;�o�u��#���\������TGI�����M�ef��L�m�����j@hz���|
z��,��{�2s4o@�G\�.��O��/�z�6���]-�����~s��;mQx��Jx,�l^o�8�kW�dx�l9�����5�/=���+��;q<�������j��k$�&>��8?4��^Qu���u��Pm����I�L<�:x�G}Sٷ&f���&�[���%�Z��,���;GL܇��[�lVs�Ư%V ���2H��1�����|����
X�۞;B�f���3b�2��V6���M'�w�+)4�>��j6+BI��pE[Wex$F-ɜ�����RN�ۤ��9\�œv����jk���ާ��#U�Z���EB9��1d��^�چ湟&�t�oJ:Z[�0�@Qua��U|w:���<R��ܘ�=��fU�J%�d[|~?
9:���6mk]"��O�#J���fQ���ݜ,��Pۊ1>� ��R�����$]���1ǳ��\��4�t���'�7�Ԉ ���n �)�J��1�46X+޼8K̨��*��m���H�0�?�
���ϴ����&A�S�.�m��?ȳ��|��H����9�iP��?�6u�4����^���@�
]��
���ò��mcd�@�f�u�+����������OG�sH<PM��E�"�-�.!1�ֲ�dH|��Z�xW�:X����Hz���^�c=�V����Rӊ+���f�/n�E���g�vE��Y���%Ok=�L�R}�M_Da���s�FH*Aiu'�(����7�j
�����,�4���
7PM��TN�Њ���劌E���>P�z�*��T.ϧ�&�c�J�iAj��	��hښ�����.���)��?�(�t8�<��b��F�$?u�[�zVc�k��A���N��e���0�W�cb�e��##��m�ր��߫l�a�s$�	(�k���W�ytRU��G�Z_M�U�Y�lEANX)6���Z7�:�֬!)E�P"�*��hNa.�l��^���(��<��~�ӱ+���Z{%���[\��z��*^����@9�b�ٙ�8>��9���Qc����BLs��Pծw���j1n0�Üv&E�t���x{�>4a�S��I�	�M[�X�3&��
HS x���.�zϗ���?�&�3<D�C���De��@�T�8Ǩ&�nI���yb�=����Z��O;6��_�������� ��N��ؽf�7㞱]5�,���+Kv��=jB��O@0�^f.��ӈ?�n��I�i'2���9���rg�5�Z�@�f��Ƒ��'��h�B~�ϣ9pV;����w?�mk}�U�	�JU�?��ھ���e����&�ƚ��-�����W;]ja ��Ns5�%R�m��q��!f�ڣ��؃R?/1R��Y��K =Hhp�[�<�O�s����)��l;��=-"��D����UML�����y�:��frͻ�ܛ8x�1�Z�Ɓ �1�BVzz��~�3}��c�����w��__\61�#�&hUq�	�>�BDj���������5�O�];<���k1P�W��I%��+،���{�	Y�Ű��\]���n�X�!�=��65z�a0P��H���C�l��
D��w�h��5;�$� :�0�O݄�0�.h� ]7'��y3D��M]�[AY�EQV	�댍W�̭�� �~���A�����:��{95��k�V�����x;��Ï{�.e���ڬ�5��;]����Kn�[x+�~Ф;p#�<�R
yw��;'�����B����Zm��������tOÌ���.?8w��e�"�`���)�,��Q���0%�͙�I�R�O�́�@(Lb�VQ.��n�Y�wv��+w�Q���<�%:�rC<˪u��H���.�<}����N'L�TJ�8�V@p98\s�_����aO��;6q��7۫�V�X�p�E/x3GݞY f7�$�b[����@����}\
{�[z,��6m�����M9�DDP�V|4/�1>c��X6�Ue�ڞ�n���Y��=���)�(E�ԭ��4��F���c���@	t�I:��ͩM4	�)�5c+x�٭*b(%l�)��܃�k��&;��Q�>5U����<?��c�bx�H��&K*��Q��d�<E��qPR�J�8�Zl�'���cZ\A��r�A�	�9�*mp�o�R=Ins%݀���7���C����W�(�R�Z��YsS4��R��b���{�ϼ���a(�M"oh)������o�g&�J�S {�͈I��K����0�i�� ���U�>ZmV�����^��xȨu����`�OK�:���0<��Mʩ�2rA
2<\nO\���
_b_������0�h����\�H>#GS�h�㼅�}5�!�#L�iB�g�IE>��P.�܌��ҍ8���qH�H��?�ˉ�M5�]B��d�'^T�㣦&ul�I�"�b�������DA��ir�La��J�� r�H�# ��� |e��|�2w4�E��P����M	)����L�ѐ��?�k����~]�����JPC1�jN������M���f[�j����h�l��| )�(��(�C0�Ż��5��9�{�����j&��6n��,�(�^��,�6�Y���X��~�>��3��+@z��x~62��eADl���?�b�&�$�vg�Ix�)������wꓫ�w�LёX��8-��Ua�onň��6N�0�Y�J���2�&ʫk`�^3��q���띋d9�X��1 F9�)�^����%��6q2�&�1�
�m���>�V���	*�F1U��=6l����CTxvj�[��c�pz��y����=���Umi#�f�$L	8`��
m~M�c������n�]x1�Sx;e�~��n��O-U��]�m&��ֶ2s%^��Y@�otD��F �c�Q/���p,3Kѻ@�����~G��Bw�k��;��G��ō���Ojڣy2�K�c!I*=W�Җ�6J]"�ke���ZF�	Џ�>�\dQ꼦�� K�T�����Z��;��Tk'`�9����q��{DdL4<��(u
��DboST�4k�ڸ��u��I��j��]5�O��'����g�����xT�ι�17('#̴S<aǥgH��&_�.?�?����D"Q'-^=��:O�<�����6�rp�1y�8��c%�"�2HͶ@��0eb�£��ñ��M#�0��Y�Q�qCۛ�������.b9s�l��|�q���z(ç�T$9����=@^���,�Sc;����W�nr��R59�����y`u�_o��|�̹_��Dn)�͋����xd(�?A�x?p+;��g&��d� O�@��$+j�iFrqߠ��TF��;�{^���B�Z
�f�ܖnG3��{��j�l1/7�\�t�K�-�e��e�2!}�����;{� �3/VA����1�Aq�hS�����~��#W����b��AK((%�٘mDIf�F�c
���-���h�GK@�Q���Y�XO����,ك�ʡ]����tw.�Dq�}C�$s��K�hC
�l�Ck�Z�R	�Z//�\j�d�� xq7���SV�r�������8��Fw��.T��e{G��j_#�t��TLz�%�w���a���dW��?&v�OA6���lZ$�W�$T%C�
�ĺl�J/��/=ǵ����I����9d#N0�Q|� )1����7ƪ8q�l�i�I�&~�4lQ#_��3�m����*���J�W��S͸ �1v�tԸh�}��>Dk���^���=L�ҩ?#�'�;��!	O���DǓ���ZW����<eM����U�?=��.Qb��3�b\�LR�xk�d��i~g����
�<F�����K�c_�私.����[�R?0����*,v? �z\>NR����50}���C��+�r]uD8g������n䢄P4������� w�-�NP���]�c���B"�94�����}IY�L����`#_~f��[�Iə	auA����O���-}�<��Z͌d�`���V�{nV��d�����@�Z]5->X$88��@��%M/�LbS��xg��回j���Q�c��x����;�y������9P�����_��=�`����zp��7�x5�P�\��z��4�s�}L���[�t�%,������z�hĞ�ɞw����r��AO�j-	�4
�!"cKQD)����ҿ����S���/U��ܾק~�H�P�c IQ��g�7B��q�B ��ʻ����u�@%2�4kKbj�-���5\k���X��?��}B�B��?����%ߏ���l"��þ׷T�{�c��e0��~�,<��^4���E�"g_�2����U�3`?E��JE1�a"�
�1Eq��lX�οg�v���yQ�j� ��8�p�#��>c�!K�����m���t�V<˦�|u ҟ�����m�l��
B���	���ښrl?P��Z��c2���
�O� v
�sZh���V��o���a�s �����N���f&\_ۂ�}2n�Y�ҝ�ã�7�^�S�{��{-�q���C��D�Tb��7q��nj���U�$����헯ή�:=���¤m�j�K��∆��"eL�$�ƒ�@�`��zu���d�mG>	v���W_6�ڨ���Qb��fKY�����w�i��6�x�v�J��\�gD��Q���O���Q�O�-�����_T}��0��6C��e.ʅ�y��'�J�U��9�:���ߞ�ݠ/�� Qj����
�����>�'��u��G�|�Q�$���{!&+,�T��GWL}�`�\�?|�05�q��.�̤-�R�MC Or!7G�X�DO���^�h�R+-EM̭?�V�m�V�_�bx_O^k�����.곷�	�]�/���i{)�R��t0��R���]/���	vL!�C9Y�լN(4��n�����-����0�VK d�z�5��n��b��ى��=H��]U��1f�཮��b�>���]�l��Z�ph6;S�֒?�8b�H��ֽ��L�GڑA�%*�3������c%2,P�c��ɻ�J�b��j5c��w�2I4")? `���v�=����S����y#SN"�Q*9�xO��S�E�O��+rw[�O���y���av���!eIPvh����M�t�~�+��? ��{�k�J�y/�0�{�����x�? �n�y�,q�u��5AS�\ר�Y�C��lL �y]yC��¸g�'��v��9�VBʾ����Ӭ�o9zȨuv�U��J�`����d���?�Pu��m��V�~4������c�Z���jN^�`^M���Y�1֜�lцg��]*r�t_��	`�L�V�+�N�LݲM|��wV�p��r�t�H6mм)O�A�nu>v�v��`lA%-�<�2�����$�8O$N�.����bg5�@#�5��lK4?���'�ڪ<?���{�j�'�i�-�X1�����h�?�·�G.�S��~<0K6�r���6�n��2�K�Y�5ڶgO�f��˼[�KqmPT&����6&��	$ KsC]lK����x���qB�Z�J1[a�+�E�b	��������8�s> `z[�S�vA��������3�Gӵ���a�$U�,֙��6?���|6��|?D���)�e\�Ȥ�R�@���\`�|�sH݀�>x�m��,МB��X�//�1Ͷ�����ա���V�!�1���������8��q����� �9*���\b��ŖZ�^��H�F�Ѹ%d��,Q�?�����lK����#Q��n��L�~gYt�J��w�d7��X�I�����
���E{�ƽ1�Үʰ1�sTn�D�η�{�sT�4!��U��*7wK�9�f���bLU���W��׍�d��Y�-�c1!�g�C#�i��Ot��5���Kw��-�C��4�_.��k�`���;5�'���a��^kh�C_�����ح��?:�X�r5j6�(6�eb�qB�A�*%��5O�ʱV������8��A��P�}	���%*��	�� �$�~�n'�_5G�Igt����8���g)FB��a��K���C6'��Ey��N���h��NI����l3� a>��qf,�������{0���z$A:9�蚽�;�~��+(x��"����YQ6����T��cA�Q��&���e�}\���!��@?>�,�db|��T��쩑/������:P�����g@���$91���+��v��d4�����Rn�����;;��)]�oBe��;2�'�n���2[������ޢ���4�9G��c_2a��5�K�au��=3h���	@
W�ۜ��˪����z�@$���l_��r��a5&x�-<e�� /�uu�2 x����s'Ii~��$%E�J��м[k�~B�qj��*��e��OlX�������9~��н$5C<P�V��MI�xk������]��})XZ�b�e]F*��9VRN*{lA��b8)��1��#�.�
�ާ;7�D�#\����r�<v��ʉ	UI߼���?�T�n��{���)1xo4<=�)�2n���g;�M��-�A�F��]Z�N����jc~�P?mU�˧��O+9,/ĺ��B%��F�ŵ��q����Pأf���f������)���4X�5��$�y��6�^���)�N�`��X&$!�.��� Ki�U7�-�)) A��!�x�3�M���]��=)���C0���\���!��W�4l=�����]X�g�&EY��=m�;D==��b+7n_'�6GWWJ�FzY��oVB���	���Eж��W=�3�B}�у�%�ᵗ4R$oui}U~��}�sY���w��rŒ��D�"� �t�s#yjV���q�o���ù���
�E��}q�:m.��X;\�@�0�}EV82CG�s�$�"Jq�M5�j��J1�::j��S��Wn��I������6[�{��\���?c��$Y��Y�VY_�7'�&6`�������~��qx�x��e~R#��]�!=#� �ĦV�_K�X;��c/Ny�~h�Nr��C���?�Z�B��>sQ&@ �J���un��'b0�������1������H�|�(�w;�1z��x|%�U�K������x��;s�
�d��R
���hc?z�,{���ǵ����e�m��X1B (vw�T4
��~
`^lj�Q�N�A=/h�������L@�[j����;Y�o;�"4�����4�����:F2d�k����cd(�̛�U��4y�`��Q��u1��bVO�F�	=�������v�&Y��!�dN����i2��2��6�aE1pA%MB��B[ԭ?�k~��m�o��f������L%CIp6#�_�=ymM��A~��'�����o5шoX�ǐ��� �b=�ms���)�'�rN�c�^�L`�iVPNj�A�b�펣"�2�-�}7IX�g�0�@f.��0qZ驮qe�J���3�C��#����0	n�lm�C�u��%�ZLX��@�y��}��j���lbrt,嗉!�օt��|(������ˠi]K�S����P�A�v�V�	�P�������UC*��L6��x����-�8V��2���U�v�3�HcqE��������S�C�g��h�(�J�󥃈���:���G�\kw�ܽ���M:V6֍���V�y_�dAv��� �wBp}w�Rӄ�������JR��9*�kֆ�r��ŲO_��D��ت�B͘�ߟ��e������0�[�=�Bq���ε��P���3�'#w���`�l��Bw
�����I��3�czC��W�_��^�l�?�	���ŽJ�+��3 �w��+>��@�5M�d�3�m��_�B�4l���d8&�!�HO^%a�;] <�uޗ���vj�B�:#y�r)��I	�S8����D����‫�m^}7����v�%M�^u
�'8כ�:Kꣿa��:{5�g�B)r ;vF��r�=
���x�;9�%:`mO�� $���$n�=6���@��H�� o��H�ܨ��� �D3cjEF�.���w}^	r"n��s�?:��"�+����������ƨ�n��'�:Ŗ<7�[7���+��w�B��p�g�6������������]5o�q���k�TG2ȯ��3I<!o�*���k���E�D�ey�m����.Y����)�2N!�l�p�y�qsu��W
�'n�]t��2���N����4�Eگ�@���t�>e?�nHo�)x��+����6$��}n3�ao���X�ņk��̵$4b��S@��	�L���Ĥƨ��b�,*��U�cj��%i��v��/
R����]�濙kN�o|ʰS#k�g<�x��Ór͓&�	��g+L��)ok}�a�_g�N9�J8����ov2�%6��6oP� z�J�M�G����P�r��$���g�7A�b/�a���"��G!���U��w3İ�@����d6��{��r�
Sg\dP	e�9g��e���v��fX� :��;其������N�P��j�q�~f�U'o���Wg"�`���3��2�eҘɧ*{2��!`A}�$f��Z#���<&��k��Mi`��\kU8'�������:�p���D+���B�^�w�c�`�� �MG��)p³�&�����|<Klv-��\>��b�����2>��V��d�Sl��/6�R_�uf���w�b����R����J�#o≵T��"IU�}�5������Õ�5q}�'hrIt
@���Q�k�ӑ�lՆ��(n�j� �=�/^É�|i�w@Q��u��P�Р?Ђ1	����=d�����unƌ�&�h[CC�ܱb������n'G�<S��;�tM1�j�A��@:xfSw��?��@d��/�t�H�����r!YGUa�B�0d�A�v1���7�G*#���YV��{c<Е7x�TS+7�	���G�3��-8��wDW�G�vWh�h�����C��iWd��i���	�55=�d	�9gZb�R�m�/A]�0[t�缠�����@\ݐ-��ȣ��G�'��$�J��4���H�Be0�C��U�yTv�Fs���A��b+��IT� ���	�%ܡh)7_�͂|X��~]\_���I�|v�`t�����y�]�#s�şK<��
���b�T�~5�KnU�I�o3y��> D�)3M���Lҙ4)�� ��>�m���z:����.KH<���T���:���j4��eX�Y/�y<<R��S���`��L�;Q�@=��Ge�F%K2Jy^C��_��|Q`[XV�1w�p"���+A���FqZ�~�2$���G�%y�F[�oj�H�К���KDjU��4����P�tv�g�E��`8�1�zr7�ä����z�8�aZ#�.}�7��Az�YJ\��koo�8��td箼�(%[�Q޼9��bt�ߨ+��!�YQ2�tý�U��q��~��ɗ"%����A[�&N�_f��)t:6&�� pQ,��{+�����I<G��E(��J.4Ѓ�f�}[�����O����?�fg�m������S�=�����\�'-�+�
O)�@�m�;������$WgOl���Et�GR���6}9��R��I�XH�t�%7A��2�s�}C3�_3���$N�SB��vX�H>e��!���{��v���֝�Q<*���n���)����!����[�J�|B$�_mC�c>���X�K�s�=���
׮?v5\�bo�����9@���ﳇ��}R���z��܍?j�L]���?R:��H�!�W�ЬL3mp�|�F�w�2#͖�ot}C������� F�y��+OI14�٥Y�Uɘ�Z�bIl�_�Q�_7�AEnA1xx"��f0�C�Gi�*>:���8ǋ��mN�n|�t&� Ǣ�+���QH�Ǻ�5_0�J�G[�Ob�s?D��"b?�w�Ѷ��js��pȧ�.Y?;�H�#���)�'E��b�^�&�_�.Ʈr�G��\!*�(N�pn���R��!��5o@G�V�ګTL�����k��/�%����\�v��߇�n	�ւ��0�@MמV2����栤>\~�Kk�L��#u��o+�=vv��䳫i/�/����d�<�|�ʓ^m�i�]�?�+���.��F�F9��,�x�ƞ���z��|.�E��(Մiv��b����Ф��뫗JM��	!^�C~�:���
ٙ$YqV��\hy�dFI BzX����<^w���5ZQԠBKd[��Pաj�:3�`�̱�c@��j���\��RWŐ�Pƫ���׍\�r���L��+��;}�N�q�o:<p�����[.�"�q6�z�bP]O���Gô����3@�L1�izǳ����fb��׊w' ��������b3@%)�kղݥ�f�S �H�������Ӓ qXf���F�g$�x�e�p�o�Ϥ/S�Una�;Qc�Y�T�Ov�0��\Fg��)KC�xU@��e�1��|��a�'�G��Q�,%ev��w�����fs��b�EI�+�ŀ���:$����,�)zX)TQ�Ϊ��XP�����x�(��h����'�;r>�5�'\�X��1��7	y�3������$
C� �ճkW��F�#��]��y�oag�e|�V�J�(�����!�h�3S�6����L�������	��ԝ1�g�+���3c"�ʼ���>�!�2���k���~QY�_ :��~��p�L?�)h��!J�ૃ�o���1�V`�逸��I�PyB����H�hJD˿tl�����B�x~ٻ��AH�PL��tX<�v{9!WR��0�Dޮ��0J!���Fi^)�M��)Q�(�L���T�W츷Jw�������N�5%�LcN-h�d�e�T���ɫ4L�*d[�%����}���	k�������)��5�*���k��rN���Y��eѯ��i��T��#��ț86?���{?�'���1�#x�d�穙�����v
X������WDA�e�Y,�	xܘR1�*=�3?�8Vdɸ~!1�O�.ߓ����LP�3*��3��q\i����鹼�de4�yt�k�����ђm�0��	�n�k��S �i���M��V��>�v8B�!2q�tV,|'�9��ʘ�M�w��/���Qv+�- MOuNw��EX�P�j(a����������&�hU���>}D��뚉�^4BR�+���( Ǧ�T�p:l9$f��������ы��/�DTp������傍������M1��9M�+�Sf��ņ�"y�}����o�Y��)�i��W��cTP@�c��OJ=M�� 'N$|��p_Kn��z9��Y�t7��Λd;����M���ƀsV��PI�J̏��3x2��ѣB�����v��ӼaU8K)�`���_ms9b��(����
��9G�5|���~���Tj.�[��RØ���{_���=d�+;̫��ۯ\3���(4o�������h��&���������ҍc��1޽1�0b�$Z�������*~�f�A��{p0Mh��E����a8������m۩�z�P����m<��	��4��1D�6m�#>ě�<F^��L��!�Ԛ=�w�#��b�t�n���b�(���f��>���eu��s�&1e,أE�'�X��ZP�����&���r��ʛ��fy����-�v� Ұp��|V���=�½�Xf�%��9�d>JEě��$�����T����i�5fʧ����G
�0������`�޾�����`��6������}B��b¥��aH�������]̎L�s�q��;�0J� 3�~S�^nJ�����ڴn��~;��g�������ďi��Bbc&��`fZ�-k����[鹗Q�/3$A��%/��	����1�"W����ف�Y�> �WS=����)��r p�Ҟ��8y�j`"���&�BU�3����/��UI�m靫�{v7���W�CH(���'�y�V�����"4$�5��L�0-�$O��@�N5����k*�q�?��61��>=��$���2*��wP�\�,Κ/�B�1�msX�DF9����i�;
J���z���.k���O-�wB-#J�P�y�����䧵P����E�!�����(���S��eW%r�J^My��Ź�t�Eۺ]�C���Z���=*�L'�a`Y5���i�@���4����:w�V�ӷ��_S����|�x��)O��:��g�������;���CR���f�Z ͕�ASd��~��%�ZnSs�U0C=]b 5d�ߴv��-ޏ�wXF)މ��z?�sw �6����n�%���]�I{�8�y$�]����t(O����Y�T��(�/��#�x�K�Փ_pj\�h�(Lw�I`=����YbV���r�.��\��4��vC��ټ�w�)5]�oڵ���  w�qXWW�x�-�}<1�ޕaj��8�O�P� �s������3e�Y����g��\��C�',|�`P*p�j?W�DT���T�F��x�䇭�N��sS��vt�e�
4ba@���V��'�����Q?�Ǘ!�WT�R���q�`0��2�gaP�?����}�U�����^�P��1m`�rk�E9��K�f�|�t��y	07O���5P��YۦW�r;�����Zӫ�Ec���k���i��\憦��3���W��ª�؍������Xz_\�[�G]\D�&�k�t6m�][H��W�hv<Q��	!b���>�a���pH/�G���:R���z���Н�\n~��L����ѳ���?���޵�yv�Dn�6U���k�<�j'���=��￘E7����cBJ�贪?Hc��|B[=u�xIA�/�b���Yfk�jՈBrL~i:����%j��.0�Cr�WT��TpՄ�}��|�Ï8�1��'���o��P
7��ZA�
5a��!@Q��&sE�W$�
3���WR����������G1�'�]�B��=�0��Enm�����]�/k��Ec ���xId�m��LP�N����_:�0����2�9�.�k{}p-�X�Hq��p��L_��/��\��t{��������?\�����5.x熝��EӞ1��~�'��w�qX�]����5�lɄ� �WЌQ��k�Z:���cD�<�F�DjDO�������[��4���M���n��Fc���מ��TfqrM��2�`o���}�&\�I�oAG:c��a�8_1p���#f�F�^���Z�O�r@_8��~��1 ��g�������L9	�A!`]/�jI	O�mkC�~�sqq���EE6��l��_$���g ͧx��D"7zNu��a� pW�@q*	f��L|D���N�B3
�B��-<�t���
au�����s`Q{GI��t�:8���T�tO����[/�c�����{*S;������M�}��=��[�B�Qq9h�cW��D�"�������dM�,�{�K�]q�;����v������ග6�xD�Pv�����J��f4<\z���h�T�DA�\���n�x�u��a";
Mk))��F.O��є�������D����>t���@p n7��ԟ�w�C"�v���og��������M,E�_4�C��s�H�3I���(�gn��X�?e�L�,|�x8���"Ó�(1�-���2��A~�[�J�H�s�*���9Za��A�౤�S';�����ƨ.�A�Í� ib�ҭ��
���"R�nu�h��1���ه����#6mw�ZX۳3��ҫ5��v�z �n�߅	m�V�:�������٧�	r|�$�W���+���;��1���h�8v�.�1��t1x	��ޙ���i�ōOU�}�a�m�]i�e���&*���z
آTA�Z@A��Rv�
�ԌD��W)��h[Yv�䀴Έ5Q#�A�(sҵ����u�0 ���O��s�3��r�q�R��,�H�CRU�;d�����p�����'��l�0��Lhmq�������H J��O�i&4�T�m�B��<�0�?���ka��mK���~��T�L�2I��D�%`�1�����@�0�T�g5z�I�<��(B���p9e�;Tm%�A������X��ܸ�=O�Z0�`7����Q��^�������$낀�=�̛��?������L~J�N/�6��h��G�7�%���eµZ������;�,��s2��+�YV:[n4V�����7}S�P�<\)h��ۦҽ�f����{�8O(תD^H.	s�m���{���#%��!��nImS3�$�z;/E��}�� �ju�#>�`�[>�q@r>���S%W(�nڨo-�tb�[c�-`|4 |i�
;�n��<aà��_Z�Xs�2�3i�]��*l ��j*�K�������u�%�iG�*:�7J��KAAw+(tàE>��B�W#,�Ս��? ���qO�D��O1���ʍ�ݞ!��'ݸPz�,%��S�oY��1����z�'��Ϭ3b���u^�����T�[!���=�мX�$�gm�FO;�@�L��-��	̯��ڃ��,��R��!9ɥ�q:A���H�86�+�Atz�7*��a�gzzdHoJܚ} J��a�=m��bA[ 1Љ�=�:i7���e'�(��c�Ѥ�γ�0�9Y�8�'���z����HB�p�����a�E��:����%�;S����mu��s��֫�Sw�0�"��J'i�nY",q�7=R�����l�F�ᘷ�jt%�?b���m��`���5A`r3u�P*�#�*r�z毐��1P ~��vu�D�ןRN�h`�@ߣY���s�V�������ȝ�?c��f7��#&w�0<�Y�lT�q�qϒ�68O���v
�;.�پe�G�/�7���,#�������-I�G4��jd%6�*!e���Eʍ�6Ld�V�W��֣��nB*&&�ͩo�ŃV��Ol0m(���hf��{���
P��S=qu��(�%EkGk�-��X��6ly�W�3�rN)4k�WHt��ð_e\���WdMM���"V�70w9��Nw���HǼ�k��1��g*���2Џ�#8�M�x����z�	V�m���/}+	m�؄_S�����v�R�KO�c6Sǟ���C�~��i�� �$�XuJmA<�^F��K�Lʏ����i���k�"�Ѿ�%��i��� ]�X@g�
��4���"qE-��0+B��]At�𻨠��fK,�NE��9���q
�Ҟdz�㌗Ye�(�/f85��j��5���)6~���^-X�=b��C��G>�SX\�v��.����S��?�F��f���/O��k_c#�̻@	]���<r�%Q �@pl�M���;)4sA|5k|&T#FT�ڄtT�})3��o�8Cl&h7��$��������W�/�:�W/�vR�H��(1Z� �q�a��b����̂"��# �7>`T��պ<��1'�k�Y��'�8C�U	��N���J�%8'嬨Yhpd�C�.��xq�6g��Ͷ�R}q�e;_wb^u� 䬽��Wۮ�K��!�˞NH� go4B����X P�^L_r��f�J���F�������|r�>���N��P��޶E
��"��mu�yI�~��qn1z�*�C���0��:]^>�?�|Q�H9{�	�4�U4��X�1��e�� �;m�J�~"f�F���!�u36�9q��U��`�g�7*:o��6�d��k�K��&��?������N�E����ng�4_c���Pe~X����O���Omu3nP%}g.�x-�K�6�r��.d`��kN-7����K�h�!Z5�a�T_�˴��z:=�nBsP;E֞�>���4S6`/��x΍�9�Nn'w�;L/��#~�a�JFx�yJ���8��(�4�� ;C6dF3Zx< ��T���朱�e������Ҩt(�Wr�a��IM�o�&Њ��>B�}m��Ltӡ
*����㇥Vnq�!��8�L|���/(��xy�kǡ�6 ��}Z������1%�y��w��_�����S�]+4J~k϶�wކB獄V1 �I{qr�T_�PBx�5.K�V�/�L^�� �Ҙ�Yn���o�>8�e_�[>�4�-ď����K�%�kUH�1��G��ճh��ޕtQ��׊�3d�K[�~�eU>Tp���̍e��ͅ�y�0,ڵv�
�XB�� �'+^]�K�������e�4)Sͫ��ʏ�#�����q�z@��Sw,s�=�ŀ�����IUZ�����ɠz��U���rL��ű�|R4����&�
��2��K;��J}�.EK��u5+%eY�m�قHm��}�Ό}�:��6�!Sr�^��TBMv:���^���[�f�GDC�m� s"���G[]I ����URm!�-�>O�M.������:���
��>��$����>��0� 
mڲ)�.�չ�l����$VGƋ;V+�~W�����Yq��̀{��Խ;����r�K�f��&P� �_���i�$�P*�6v�g����S��K �lG$m`p�oKra���F���0�0���r��T c�m�f���J�����&v��c����f	��U���i��=�F�v���Cj��������� �{5�M>��+!'��Jѡ%G�;jJ����^�U�9a����՘��5��j�o)��Ǜ����Ӫ�M�p�we��'c�!��&q���yT����*{,��w��a=F�c��79	:I _b7G��uF�����j�����/Ώ�Aǌ��8y()*=�q��Qw$�s�;���# �pl�ړ���f|>1+y,���ٲ���ͳ|}U����S�\�;�QU���%��<W�i�{��5A7��}!��ː�T���Q
�{���_��9G]4�h��M��R�¥F9"���{s�ͩ�K��.����xpL/j���a�eG8_��0�#��_KfB`�s�/&�Pp�0�����L���R�0dϳ!�կe�1eB�csYUK�9�Hh_��͝�̾�؂�@������BMH ���5
`e�>t\��z�H�ڽ$���2�3&�Ʃ�N��^U�j�7Cu6\�[�-nԬ�G�Ùo��<�G�$��~��#�v�ߏC�;p�i$=^��p?��5���Opԥ��b��B�bR��}�Ϥ��v��J�G4�$�&�����b@�y ߚ���ĹF�f�My��x��ZZ�!7i�
���%��{�C�Z8k����\Gؾ�!ӿ
d�UM;�EyP&gX�]`j��̱�*�<�,~��4w�A�l�ГC��
���Z�h����[�Oh�����L�k6;�x��I�٥{P*g=� ��x0+�/��a;��|憕�?_;.����Ψ�$��BS���Ջʵ��o-��c�� 5~w�2<��M _3ˌ�r�.a�W��ĳE7���(>�ؓh�Z�� ��c��r<�L>w��V����]F���&AS*.�����>�Hɨ�"�����G/�*p���\YE[xvr�#Sw#���.��^�ȼ�T<1�����S�_���G��w��%:�YZX����|��'X/�䯘��h�n�S��-5=t�gg=T%�t������~�(~l�Z��x�-�4���Y��`h\ ����}:����������\x2A��I�p������ƺ��
�k�	�%)�-��W�w������H�$-��Y��p�\��Qn9�ĤϘ4������p��;��z8�����mHl*�{or#���r���k�2������{��M���n��f?�&j���Φ����jR��RA��'�\d�%q}�Ƣ9�����?�sN��^��m\Ƌ�T]ץ���g�6��G���Ҽeef�/�$J<2�)X@�O�8P8�;0��N�u�]�C � � @m�W�C�*���&�x��0�1*o��t��a�,T�̏*�J�[!˭7��+�e0������c��hәj�,�*%GjLd惡&���ˣ���y����B�j3KT�mM��]�2U��m�.��o�:�Ӵ����&���jey��qK_մo��������c�V�V��$�}����U7r��}x�PmA�V�^_��`��YKe��Y����D���^V����#�J(��6�Kk$��n(�ߚ�73M���&1�"%v��׉�I4 �%��#�#��`�ރ�g��ί���}V�<e]߿��k���T����[J�,��˵@ٔ�׎vr@U
xk�ܤ��U��2eS�dW'1Mɵ�dw��
�/~O)�Ɍ��$�a��&���o?���p�cK�ѡ���<�ʯ �o�$��Y�TD�L�c�SR��PZ�����џ-�xߢ<����6�|���>��]N�V�DA��A���f��,](��?�~+�]yޙ`f�B��Ԝ�R�`���u
ǘ>����;HoB#�5w�[�Bo��}Q��X����?٩'�+N�+4Y!�n�.�b+��3(�Eꘝ���s�ya��V�vCC{97�
w��hu�KZYX�#�2�����~�����-����g��k�ҏ����b"3�sq��0�ou��|0��iD�M�գ��Y]R���N�B;�����������}PY�{�R���'�)dR�c�t��=q���߹VwR��2�b�u�H�!6ȝ$t�y&Ո�l͖�S<g"HF��i�N����i`�ϒ��-�auk��i��m�24�)v ���폋9�Բ7���ٚg���6��Z�W�ԁ.{E��s$�]Qm��qH !�%�l3X���B�k1�%�5�
�E�<P�v�x�s;8��(�X�z>x��h\�������-�4?%����lgt]2�ޝ+����R4D�|����1�Lr�Q�'P��Wb�o'��#��4|�T��;1�yd�����Z����6\*S%}�jQ�OsS���o:��.)�a3|��!�-�B�E�����q-�U3;h]A���7)T�R���k!��P#�����n�8g�I�����H"�/���de	J����|�Q����1q��= ������X��-�15��Q�JC���D����1u�*˾BW��L�G�H�V����{L�y
~��0̩# �l�.E��U�6�n�<a�Q|n�!�|�|zI��}Ԣ?lƚ��T�ʲ'ȭX�`(�.�w��p튉��[�P�v.��쏍4���2�s��d0��5:Z�W�f(�������42��*->]kv�Z�4�c'�u����sw���9�r����J��W��e�V�xgZ,X��[����`����?��~Rd�6�f�W+����X�4�Y,��2�g-vԀe'�;�\V��.W[�זׂI���8�� ��T�ڭ1�ȫv���Y�����֬�G�D��������h�"�b��9�s�"�0~��5a|�ыG�J�����(�,���{nTM��5B3��w)Oov��3����|3��*0t�.��ʋ���[2����9��f'��������$�撥�7�C[v��.�w(�".��9f�����׼B����QT$a�=�AW�0$^-��w���*�

>,�Lq��yL����M5�;�X�j�0e�o���Wj�Ƹ��2h�Q;js	�!!�H3iMM�����f��|���<�ݔ��6��\���[�,R48�@xH$(��,���6O�(ʆ�����r�Kv�֗�dR8�G�z5u�`9:Hga�Ժ�fYN����%����X, �Z��Ty�w>�­��cɧ�<�d%�5
��.VW�P3��=����+�D_"�ь��Q����,�K�V�tN�.��Ne��Iw
������Y���-�rXNI����!����|w��!c����]�G��T�����z��6����p&�z��_�Pș��Z���@��f�*�,���A̞w�-��
��mF�,���?cl�'ʦqA�x���2C�z�%5Oc�,�H/��Nv7<Ӹ�o�bJi5��I2�r��UrB)FG/��_���2KߍW/�����]@Vi_C
�!W�b7X1�{���[�*;ո��{ae��K�[���~򌳷H5O3\�^���������SZ�9�u�֚��n��1�i|��J{�e���Tb�q�}�=)an�bM��1蹤��
���ax��͚�H���Γ �0�۽=e���v�q��	97.ɲ�Dߩ�en3I.R�>EAq�k]�4�5'{mV*g%(Ó
J�p~�wz�y�aӮ�|�̔f�,�w}�ˀYB Q�
R�{Y,Xc���Ra4�hN4&�ݴ��-�g3?H�8\n% tP��i�(jl�GL2.Y��	<n�@���Y(��*	�ʥ�[�/x���	6�4�����)��6���6�%�`+!�a��~(d��'�%uF	8�y?[�����{�j�68��"jԕr�Ǐj�ޛ�X����$zOV'�3^���U���/�J���ήj ;ɚ�p��S�.��?�'n��̂�4���i����x�!q���)�e����L%���	Ⱦ���£<B�_O
����mOH���b�����!`�C]����A�ɬ�D���M�$�������Gs+j)�����k��j�qt��vE�-?�5��3,�{�9��{Zx�n39cl�xk��K��Q)��%�<�'�~jՌL/pʧ�6Y��(D���5jt�`BT��cs:�!���$�]i/���yr��'\Ү��H,���� �
C�m2p�3�Zk�-h ��]��Ƅ�*�ٲ:�7fv��4��7lV*�~�J@:����<����^�S�����Y��J	�Ƀ��o����/�צa�X]#�6g�4T��N�@!p'H��:��?�L�G���e��Xm=`�Қ���]��HL�-I�p1�5o7��;��9hr۹/^��wK� ���[~�^���h�'�*~�,�{ܛE��=�iU2�79>$��
���?fюI6Of*q����[?�JD����"c�͍� ��=ꆢgi�e��%g^����~�m��S����7��[�F`ݞGYuzJ ��&,$ �Yc�#)!~����q0^��Z��R	ݒ�^�˻�<q������e4���£P�a�[��%~q#	��MF�U��n�~o�"�h�8�'R�b�rA确�2�_�3;y�d�1����i���;��p��Ng�WU�K!�=	���d������+�%z]I{L�u������̉)n��j�l_ �i��ߏ���2�d.�{`���7�!��^�6]�Gꌼ/�O�R�ڛ����l��B��x_���8��L� qz�ǽ�޹x��A5qY<{�.�6n��u��_cO��Ǫ/Gyt���o�-oZd����e�ױLM,�zn@���E&�!e��}�se�_�G�u8�yѵ�8��x�,OP+��Re �h��*E8D�eQn��7i��C�9��\y�6Y
��l�G�=��R"7�{���)��ޠ؟1��[�ݚ���h��������wA9��Y��R����qD�f�_1k2��Խ
��@ \�.�m�v'����/ۮ���p�n�[ہ�*���p�d9�C���Q��Ձm�������X8�DwoW��qt�ۂ�cj@|�E[�,z	�Oh&�k���"cOVt�z�����R�BUY�Rw�_qe 	�ZǊґѬ�� 5����` 7�$���n]6�FN��Z=3���S��JQ�������N���YA��n�50����%�7�k`�qnu.M��lN��4o3��s�p� ����Ϝ<Aj1��l��T[#$�z����Y�����������r�_i�#0��փ�� f��` ���n7v|�<�H�T6c|4���q"��!~,U��zY�6�tRaVo�������(K�!C���u���i�}��bϓ3D���3C��<xۇ�e�@� �p䤊�D�,�.�컷���e\լeEG/h1��H��R&�8�Ȓ�-��7��~j�M_"�|UL�>�6����Y���:�FՋ/Rʩm<�dL> �<>�+.�b��B��4<��4���,�2�[�BO���cRva	�-�݁O�xl{�ʝ�^Ā����ai�}p �KNQ�ޞCR+�"av�����c�;�Af{*�f���!%R����*N'��4숬�5&��xz�RQ?���|��M^ևô�j���Nm:c�P�̚L}	1��M��H�ޮ.}�O&��^D���\U�"P��#d�03�.)~��+�CWj+�{�T�h���B*��m	�Q�mgT�� ":bٞE�3�4�o����h)��@(��g�~|����m
r��˕rn��#��&������Fί�t�d�h!0Lʒ`���nK�Ҙ���:���%�[�Y����\܏8��tf--(FSgk����w�P.��$�����' ïohvgs��@�[O��!3�.6R0��L-����'|�&�i��q�B
)�����U����Y6��זm��?��3��"����{�GKܶ%������\�[Q�V�t� J������T�}E�݃��"�ˎ��x6I����ᚴtI�W�cFBH�4�VLU�ǾV :�gf�����j8��4��s�6q���_l����OM3;ѿFC�x_����s{َKGL�c(���"����p��0��������F3NCN��C2.Jn��_� ����	����W��
�L=�%�G�(n֋�'_�8���7�O+\��7%I|Fj�'���_)�J�b%�o�S��[;~N:� ��p��ۀ���y�7�@B�k�|pF蠜�z��.?����>o젌�o�P�3:��
�X��N�F��HyU� ��+�������-�͝����~��M���I�is�[��B.�#t�}�����U �+eLO�kU�-!���z=�&;.1�(��jϐ�-�P�s�a�G?}�1�o���a�&5�bt5�����.������hx8�܆ꀧ�?K��C��@��h��H2�J$�����vs�7|�[�X���,���Z�\�Q��e{��$� �n�6���%bW�T����S�oC���u�O�t�i}ฬR�����q����#Bzf��$ѩ�&��G�D ���n�]4�6)�[�d�Ը������RC!��f"���Hk���eB�k}�tէn������`a~o������>��4�W�W2��$Td~,N�,�$y��Xs :�z��
�A�l-�psGm��7��"n�QIWǜ�UE2#t�`_yO�#���Z��c�̓�V]��{y��^`:�aWK�ɣ�#�l�d����H��F`ݐ�2��^;����:;�}��Xqj�r��0fb'�;{8䅛�%b�����[��,%w�Z-ޑ��5�6� %��ӽ19z,�Q+�Q���gj���JO��tDr�}��Wc�J����?-��C��HZ.`E����@���3�vN��K��-�K�����v;B;�����4�c;�4���8jgTb3�fE*�-�QQ�����+�ŏ����F�^�orQvK*��Q%po�k���q^�����C+.�r�B3�h5됿�)q9��8��-J��Y9M�n�	�El
�%���ӥ���0yq-�=�9h��bF�N�L�K ��S�#t�բ��-~5��gZ�2��Tټ��= � ��XdH�lb��Z�]��P�B�i�M��v�9�̙����g�9yrˏ�1�[{z}P�����=�;$�Xujj��m��\��i��Q+��R�剼sЬ�N�)�g��VO�'��h���==my�f?�����cg���_v��F�J�V��N��[��ؿ����-�ڎ�����?��2���!}��)g\h�PN���Vf���O�8EV�	:�T ����t���~��F"����+��'�g!A���"˛uA������(��X�yF���n�(�pdR<N�r����S8�_n�`e��㲬j��F��]֍�՟ŉ�����/�ˉ��fW����5�Y����f޺m���n��������ۢچtK����cSpM�V�M&@���Y��o�LBT*>�N���,i���L55[�����C��b���]�M%���.����.خ���Y��I�$��s,�✲ϵ�)��D�+���̜�|4���"?-���1�mB��Xj�ҜL߷����~��X���� \�������b*O!��j_�;!%q��G�|�k��}{���W���K��Ř�V$�1�5�s_��p3d����(�J��Vv�{RM�T(6]{�Qy�N��r�^��G��[�}��Hpxf�*�
�,�v��oU��&�9��ӭ����{��JJ@�խ��,�c-FK�X�
���Z�]�(k,g�w��d*Y���̏��z�G�]�[h`��4��,Sc�Y$!�"E��\� ��y��4����]�X�T��{����8����<��c��'�� [Bg���
�I��8	���՝&ټ�4Tҧ$�M�ؿ0�x����xf�P�UozY�G�3�aX�/���+�Gы����cX�[�R0}���T��S��qLq���$FH"��w�,8���w���^�"r��m�|��?k������,��dg�|%kA�HҴ����9���i�Q{�Q6�� \�\p��f�ށ�]!H}��q�ZJ(�L3d�X!���o��K�O�NQ"��s]���uȿv?5��(��,v)P ��z) .+g��?�x��T��{$>�/�B���,i@�e���̶���Ef$v#6�Ȕ=9h�ߒ��2Zq�:?'~���'߮���c��s���'�aЦ�����2��D'r���Ѫ���K4ϕ}�ϿxI�?�Pw�g���%�ZF��79�-���&�����?=��
�K��@۰=��*a���:�q<io��|O}q�N�с�Q��X��#�+�J���C�]O|>r�yz�q���+���G5�Z? �Bq�j����~���/9ȱ���xlG��x�zj��B�u�W	\��=ct[���=mw�v?�L�Z�<������}��Պ5"��%o���{(�Ӆ��zV��D��?��h�K�gVŴ��?��c� UTY���*r���#T����J0�����m�X�GH�T�'3";��	�0����=M�fE�-��9�!"��G���d�A�=�tgYQ��"�Xe~�F��}Y��s��#,�)_)(b`����{�űq�h�x��X�f���S��Z=�sFR^�l�'$|7�"\r9�)b��8�z;�Y�EA#�� �i�uU��K����n�[���q��@��KK�~,��R?�Vl�:�!~2�34�6�9��3�b�苉BR��-������%���k���}�%q��g���z�O�����Z�i�lX���'������T��RW�x1�"�s,M�ı�G%ὃ�z|%u��%�5��F%-胻��Ԛ���_Q#u�!�ꅒ+L'�6l�'���#�#�9���y���V�)����'�����i$�G/�0n�y�|� �q�݌�9��g��,Oc�'V���85�"F�;U��f�6yF��ɞ0�MC��8�����݂!/e"�L ��0Ƚ����=o��L /�Grq�܇eGS�r�Tȗ�4֢�1�F�G����e�X������l�^15��G��B߯�Yj�����Dʆ�	��ﭩ��Qӕ��Qw�A��45�2�B��c�$�b0)Y�!L���@�9�K#e^� @T4о�xOȁ1 `	�v�T���}f�*|J�O�8�*��y=�.�W���K�9V�"�^�hr�M�����?ݒ%k��׀b��7w Q�ȆYe'��=�SA�LO�*EDF���L��r�hY!�8�J���V�����l�hN��so���\�z�c��s� �����\�B#��QMs� q�	#Ą`<F	o�&m5�X��z��m�92�+[��a}9U���G��~��Ӊ��+���C�F�b�Lt ��5��o�I��B(Iw�R.`������N@�s�STnb�������wm�"lP/���)af��ދ'y��r�#SKscvф�ךr92^� �-�:�
���^ؠ#�N�B���l�H{]\�K�eb�GYQ�,�U���g��aeJW�CO���`6�G�c�P��������!1�Q��DҭTH�p�L�J�S:�"%����� �Ɇ>J���c<���ʞ�8�{��7і<ږ}|�/ܨZ�S��\a��}G�����|�Pa�����z0g�$�6P�̛ŧ����:����]�Vlб���˯������ �5�SaD��'` �qE1t�`?���άqBM���uiڦ���$����W�zB3<zPjՀRL��BZ�S��$�x��j���7����(��nK)�@aٻ����`��|j-An�:c`
IjQgN~
��d--����e\�I�R�=�n��B�@�o���.X���g��?N{��5��k�� Q��ܾm�t���d�5Olf�|���T��s%�w��߷��C���Q͊L�@�f�Y8�겶��6����U�v7M̵k��&QɆ"27�͝i=A��X�cՈ�V��	*b����G�>����X�M��ZRfo\�uX���]�d��Q�A�JǺ8�0�c�P�闵wƈYNZ6x�O����j:�mM,fU5s �AҭƯ߶�y�q�1��h�^~l[l����G�����B�%�Ρ8LK�騅|ù�
�c�@f���L��~���lX�`:W��Rb>]S_ĵ����r���ʃ�"(l�Y)�K;rI���H�,�=��`�Q6R�S�u %�Lw���wA�&ҹR��84轣�H�V��H�hr*��l���?�<�A�hHo�oW
q����K�l��d���(�dd<A�4%�*-jJ\"K����K�	���=U����X����8Ĵn=����}���Xtw�(�md*>2ǡ+XlKX�vݷ)6���.+��Vf�0q��0�BK�[Y(�,����s�:�F^��~�]��p�{>��:��6�70�~��N��<a�x�~3?l+��W���񁾿�D[�1�Y5�O���M�d>�Ȍ��3��"��s�L�����PrltM��	
�����7*�ƍ���W\K��r�Z�����e��(4��1��&�KGz\�	"�JF1�ʚ=u�W���/?�bڒ���1�eol�����;�j�g=Z2����cl�[PD��\�KY����~�>�=���S�9���bR�E���a{�ޥ+%�"����F�Aw�4]���܅�+��J�~8@I&/?R��巀����淄��9w�	��O+a6��
���������9.�Y�J�\�.�\T��bC�KY1���pV=Y5��V��d}4��lL�y��ɮ2K`Yا�bX�zIˡGy4zw���@q5��Rl���e��B:��1�ЪY��nX?|��>�R�"̳JHJ��\���-Y/d�4���̦`:m;"NQPɫ�^Ll����eZ���~�7����Q�"9hÅQ�N��G�.A�l�F��NШ7:�$N�u��.ۢ�z�O�ط'�ѣ�9�O����ڜ0m�a��嶲���aQ���IѨ��S!CIn�k�T�Q��mB�HWqxeĚ#�B�<+��N¦FF���V3�_e��H��V X�L2�Md��7�с|J�̫��P�~G�1	��PxM����T>���I����j�d.��+"�7c4��@�5GwM΁O�)��
j�&���wT%;�1T��Q��)4'�V��qv�j���
��t���'p� �j��;W:�1:&�3����A-��'��}E�n�J[p�X櫼��w�b)\�}��i^�bLH��J��ɕ|���u��hKh�����x��KE��Z���RZ�d��}��5x�����10O$�iU�����|���w�a��-پ7/H���V���x,烘G$�6�B�t;5�.xYe���ݻo�>����0���(��Y��A\t��!���EjB)��5��*Fރ�e葬で.�ngr�r;N��~��B�9�(����1X�T�=�ޜ3�K��1���ٶz�흣�H1,��i�zbba�X�IS��D��6@L�*��0�2��䱂Ȏ�.]��q����ܯ	�#W��G�P1|����	c������lyO4Ndb�
���ܟ
a���f]��eMZ>��36;�L���:�����mX0�F�#��dE�:�b7�|U&[�)�n�g����r�ч���U'		zl�ۻ)���B��J�2����E���Q�f-�h\��=���:x�5������M�l�x�fɞ����y�S5�B-�	��(w� �58h�-�}F	e����/�H�r�=��8��n�*��HPxT�d��n�e���[?z�E���]	��d"�H�^\<�=Sa%}8�;��=!����A�zپ,t��JD ^�?��_nys)�9�U�8��]���~z�z�����E_�c:X��2�Wg���ަu-���	Q ��ʠ��]ҋ�/��9�5���2=�7�A��ͿwO)�H>Go���O�%�����y-����������g2�5΋�a!����I�br���[����"MI��í��g�01H����iq��`y�g-�aԡ�,�t�%Y[r�GJR:~b�:��T�:jҩ�R3z���W.���K?�`��ϡ������H��C��{g
��g�7n��c�̒���r���w�Ȓb�3�����yx��O(�58\�3M��yE?8$�376������c�伀�_(�wj�_.[?s�ߴR�S7��*�
��f��C	� V��q�Ӻ�b���v7�B3��sf��b��g,�^E�(��vy(�'�`'Jqo�%��8��\�n��}�&{&�����P���@�Ԫ�p����_�R"�:l�����"Aq�D�ٚ�%h�BÞ�G4sJ����-�Cܛ;h:�F}�O1Ԯ����KG9�������"c�!|Yh4��N�A��\C�����M���:��`eA��P��=_��ws������*|}8fr�9{J��������a�_���̑޸�LM\��uwLU�7��8zB-�m"$�q���{����&�D�.u٭��,��5h�^w�K�;s�;�$�zT)^����k֤zd?*ه�W�y�:CC�w�N�j�ģ�1�>h�1�#�Z D� g�Pա-�~-��k�QG0��K
�\G��`q��͙��t����C9�U�&�~}͞Xk���j��i�:kE�տ�q�?'�����B���57�2w�]�+����8����Q�pj�o�E�F�W!�h3�G,lk
�\ܗ�]�ILxбo�{@-�4sm��J�R��Y�@1�ީl�e�x�rh$�y�E1b~�zB��K<��.4��+n��?9�������U^.%�̸����={������մl1�ցL(�c�M�^bw��%"���oB�~1��7���.�'zr�ܚ��>�:vC�{�y�T<E��zbf�iQarv�C���@�0˅bR+���=�^<�g��@����-�#.�+������~�T�1�1@�3΅�χ�Hn-�(���em/?"HeJ�yVĪl���P^��Mo�2.�>������`0}���!t�j��(c���2kFL��-H�yf� >gǐ
������u�����X7%�3�b�S&u��($��70W�(���2>`�VlۂJ@J�G�V�A�w#���W`2Ee��)�--��Ő{�:�����{��� Q6�ǡ����(������X����;�nm7%Q��<��|{o8}͂��ֺ�[X�9�P���C�p1�6@��u���|oV�dga�+�m�Pb�k���^q<��>��X:o��keV�
��6��S����$�v�n�tG���c�o�xm%�7�+�G�[�|U��`uّ��N���2�2u����gchອ(N�L=�@S7���z���pX;�J��n��UU���OF�̬e%��
��v�ev��K���|��Us�8�o�0�-��/O����e��{v1����wWh��RP��\�T\��C��n��ȧ�3��R�"�G"�|[��9�[��?�eH�ثf�I�����d�\�l�aI6:{�""�������:��@���FȺ�th�h_�"�#ǳ�	�0>u�rj|L��JI����<�.gvG!#���{�n���<F��D��:�3����y<��#G�P�q�z`ǘI&1������q��Jq�vJMP�0p�v���<s��X����:�K��N�$2B�q�zf$��Z�r4$@|N�Otݑ���5�I���U��o�J�;j����ܸ ]Q�p��Nsx��&V��TBR�����L05�
��5\�e;�c �n2O�a��4�}�WP�����yjġ,V����g�)ybp���g�#( ��}6$F���(%��+k�\#SA�F��F����gt��uwG�d�{7o���xznɎ��qYT��h^��U]ڕe�w����[��^'V�z)Y���>���Y۠����>Y�,��Oڥ�+��L����^���K��!CEy!�*_������ ������YRF�O%�y�Ž<�'��C��`�O����tO������3�'6�]��訤@0����z��a��V"�!Q�N���vZ`�aa��>mݬ
�������3Q�Ul���h�͚uܻ��|�B@90�?)UQx��i�jAǬ]��0�OZ|+6�9��/��['��o�vp�������������}�!Oor�d_�ۑ\D�0�͑�{���m8^���Q��������P����DO���^�7��������gi�kB�,s�y�FV�[�#,�=�������:_��ڑ���/1�w���T/<g����������Ҥ��e��:=�?�z��c�|���, mS�aM#��5bX�ZڿUU��� �b}���	@��'�q������� ���j���UH������ٗ9�����[g��Z�o؏��@�ƆZΉs�_�	A#̟#XJʸ���ѡ1_���,�Y�������җ��c��@��0��&qL�6�M�x���4��3Xn?�~��8Y�8�;�_1�Jcc�V���F�zK�F&���s��ѣ�Q .����/���M�f7���l_9����+ĨHA��E'z���}��w:�*��ߐ�� �0��P�0J����b���1s�G����W�rY폆5�d��g�>+Mvϸ$ȇ�+g�`�\��A"�)�nz�=M|�ί^�$�=�\�p���$�@CC"�F�Q]���#�q�J-���I��$t_��՛M�/=0�>�я�� FT���S��}��OT؉�ES���P�fxK0��_R��@	I�z�ٰAH$��:/���E~�!/��%���q��1k���֊�0�C�x9�A0�[�:�(�`Md�S�f�������ZB��l�;��ld��B���g�r�[F�MǗ�\���t><����Cz�	A@�t'���|�ܙ��ю�ZU˟E����u{��!��v�j�9%b=�1��y��F��6(�F�[��A�VV,hY��,�(��tE�y�C��c��@�=�9����Aۄl�b�}a�bn���*��~��K�~a�+�����^4�
��)N�O/�d���������L�J���;`�{�N�5<�O��sK�<Dxq�T)nðÂ[g�rwzh��#&[A��6֖��F/�SI�h����X����֝��Y�M'b����`L��	~e��� ;Y������&#���$Kvv��|B砐���g$!��!c�~����M���Bk�K�:CR-�&�^�Q���_<2��o�S��!�\Y��&w#�o�"�i������ ��
Gn�&o�~�Vs������,E����"Wu?W�A3��˦��)T[L]���lo�,奭�AK�R
�Q��B���2�I?��::�2V�|5N�/��%����G����Ln.VʫF�	��A}��vM3\���&�-��Ð�85�e�GZD�� ��Z�?������U�eV��.����I�ˎ��W'���oY�I���]�+ܯ w���O�X�Gs�>��}�7��u��sZY{�l�����S"ob�a"�w��?H2��M��N��ѨU�d�ldt��:�/�y�$6�� �+Bd��ܔ[L����&ف
{x)�[7kkF�д|��#�B{5�����U*�ُ��ç��:x��#�����>���gx�e�eg�fuy�[*5��H0��*�d �>�޲t?�:���VTD ��H�"��'�L�rʐ}��h���*�N���'�^r��&p#L���{q=�t��8���Y!��a$�@N� �u��0qIU`��w�(3����yQZ��j|�01g;�N�+S�\�f������o�	�B_�E.�c�&�4�Z������G�/K~�=����m�8�QC�mY��6 _��!�f��n g~"�qD����dI=��O߲t�8���::�Vr@n�򿖴Gf���x�B�eW+��\�c��`,3��<���&	�>\}�zr�{�.��'q�
�9�����cF�سJ�e�� �zٺ����)�6�5�qM��=+�t�?�x
��cm�>$P�kC�/h�� Dɢ�q(�i*�1�:e���$�v��1�� 0U�@\z�C8��[�h���T�ex��1��9���A"���Ҹ$�5�}l�o5Es}�����a����#Y-f��z�מ�J�x�%�?))!P��fs����-gj�n,�VI����c�[�Dn�ԅ(���fЗ	�.�F�E}�&�o��r��O����1�H�.>y��ߊ@��s1ŗT͓[�\���1LZ�� #��8��xl>e��!�[9�(��\�˶���u���^�:b�f��`<����O}�����ǆ��I�1�oCҾ�K����(p.�ˀp�?�0+�,�('3�^͵��k��}V��W�U���`���bl�eǶ�s�80�ߓ?+N�CkV5�z),��� ���2�4U8��	���4�H�V���k�3SFR��p�2�7�h*E@�*:�_������/Ms����_��^�vb"Emc����3x��X>��̭l�ύ���{$��g,+�b�u��������'���^�&��&Ϭ�a�f��7VYXv�&�v _���?9=�VN/�����0	 "C�0�?����6&}�6�{
M��~/B&�Q�W���UE��n�d9�^g�s����R����b4!͑X=��f/w�z[��-�+su�� ��xd�H��Q����Nr��K�s$�{�YK��E��9;��V��aIE�$r����
���#v�o�I.����>"$7��|�ԉ�%��C\����tϧ�E�4e0C��fB���A�7}���u�Y�����j�-��vy����t$e�|�40�O�{�Uw�L�Q0�t�H��H��[��� wz�9>/�K��qĥ�6�@�-����Oo����r�?��3U�_וT���վ�4wK���X���r�m����+N9n�q����!�ŵf��Z���3���dT�aX���ve��I��ε�+B��q�h��jfô�M}31N�3���o�T�g@ߒ3t�G�n�V�y˃��<��]�ZQ�j˦=���֪ͳ�Zlϧ�R�u�̈́>���Rݰ�E�l�~|<��Y�Ԣ�cl�Ԁj��me��(q�R�f�ϥ$Cy;��U�Bʾt��W���R�swK�O�xR/m��������̾B,@
rl��R�]����Z/� �,�
[73�I�-[���i���Uo�ިnײ'^�^M�-�OQ��ݪ)���+9��D6����, /��DL�H�h%+�ޞK9\f����x.�S=�E�.�m�zI�{e"8�Ɇ"��a���g�'�\�{�y#�x�[t�-A�$�J9���|7i��2� "$k��y=�\�}g�����j��~E�R�ʿ?C'�p?��3/���mW]��T|,"�w������a#8#7�J覎�L�K%�8;���ҸV{j"�I�9��H� E3J{��x1/�;}�%��#�T�L��T	NM�2�6�	���.d�u�'���qyl����SFQ�E��l���~v��7���⠇q�pG����y5��ol~e�\KSJ���ֱAN�\�x9j�]��j�/~�iR;+��豘_:��	E���'�4�sdШ�l�s�����e����X�9J !>��OfD���8�\�Ko<��L���F�a���O"s%�!֑����+�Ҵy#L�(�$%EhA����m|pЊ�f���Y�
��$��PrQ(��!%熵R
'b��ݏ��������YּI`���͌�O����/���v%}�"�,KbF�nf�ŴI�R�k��#x���6X]4�ɸ�t�ֲ!+�ӿ����
�&De�&����͖0�vY��k?��4\�dV�`��jJ�さ�y:�Hkԋ#�c��Z��QP��{�`{Vȸ0�r��*o�����wF�h��=\6����8н�(z���F4`�<��W����'�ڇ�ΑT�v�j�*���M�dG��W3�X�ӛU��r�d ��ҳ�q�{-��B�n\��"Nw�UR79�F-ƨcm6�c���K��L� �{X�ۺ�ו����0h��՗&uQ;Q���Й��`W'j��D{�L!�� rߣ�X�2�����Z�_��Յ���l���P)�h+b҇^�6��7�N����!�����yw��Y_����zK%����%��5�.�R*`�lg�	?D��!n?Ix��!
TȀ�q
D�zjd��ʭC��U�g�Ę�q@��GyY>t��l_Ը��U�n���>��X�x��X�m�^���uΜ	?�J�)�j��h]�P�4�ı���]������������b#�g��fa=ɘ!z� -�t
�|�h
�9��`7c'.�Y?4f][��C�tmx}^/|j�A[�����)���A\@���Y?͌��|�� auϩxf�A�| �b��t��u�`�g��p+,�N^lޏ��LQ�&���Y�Q�i�4w�Sv߳��&��Fr%���c����b:�]��~n_q$D�q�)���M{��Z����v���9 ���V3�ߑ�_wF��?t�j3gs�hؐ�Y�z�E9G ���f�W�M'z���8��7�d�4<���i����u�Y�8X���P�[�Q�����t�1d}�{�WH��9������h8.5[R�2AM����+q0�g
�`�G�!��j��\Iu%�G��d�>�ј�2��ȑ�	[���	n�V,�j>�e��_�A�ރ":j��c%I^0A��\ApS@��c=����6�٘�N�'�.]�U�$� �=DM�����+��iv��*e�$�NA�Hh(�b�����ܥB	����+5^V�A�'��>�	g�<¼�p���Y�]�Ƽ�����Y�.t���=�
{ɷ��_E��I8 ��qRi�]1h��]+��\�Z��*�q���aQt,���KT����pF�_DG08#Q)���fYnbӇ�%ۄ{�c�&Qɭ�2���t��w�쿞,x�3c�j)yפ�]����ͻ�i�}�%��O�s��v����-KNktY��>��$���cmϯ���N
+`��ӿ���$U�mw��������,k�@a�4��B��C�*�+<�O�נOE��-DsU�X�{q@��+a����m�SW K�F��-���{�$��4�<�.<]0j�s��P�r1c)M[�B��H�mE*dI�8a��Rt��]�to�0�[0��i���Ӫ�v��r��<���;?lK-W����pf����%��:�j�vԆ��%y���ʆ�N:ؖ6d�-�B���b����M�zoR�m�.RY>`7W� ��ײ�� 0� �{�wN��AϏ��~�Bj0�*#z3f���������N�,�b��X>�F[��_� �%l�8h��y��`��H���	�2M{�(rC"���.�v���6+1�+�/f4�q$d.8�ev�	�5�7LKszr�,c�:�6�z���uO)vC��f�Yʆhq�貽�aj45&���xd9���lG3���:g&'
H�E*Y_�'�í�I�F�t2F��%{�9������o����-�B�����B-��p�ψ����^/�I�H#����Sw�*���bC�n��[��^'���T�z��[T�:�Q��%\�H�>Y���Z6�0�[��q�A�?�-�Y�!�`��cqז�������]���;�דּk��=E��ݿ���W�v���l��bQ�g�c_� �:��G0$�L,������[�zB�ù?cxͷD(��T@^���י[^6e�Yd�$L�RvbҰu0�E�4�� z�\�|/PJV?=~WS��O/���kl -t��f��9d<�������ל�6�Z�	D�@,_�Ľ���	��Ë�k�+�e;�Ar� ��猓Q/l��1�3�Qk�Z��,�^�f�B��p�zJ�!���}���k��'�T@��0� c�cko���ϱE�����|��q�KI=��K�#��&�����h��qzg������H���V�70%�4����vRȆ-�ʦ�G��L�g�ꙥ��lJ/9�;4;��Ǎ�Q_t��/a�%��x�Ȳ���A�.�*S;�в�PY���OJ:��:w8���o���3#��V�]A'�K�>kF`�F���5�T�M�i���j����~c �؃O�~36�O������Dh�;]d���N��͠0A._�Ⱥv�)�K+����~�8&�2x�T�n�N_M�\��t��ݴ�p)T�����1�%ݴ�m6��op��G>U$�'|<IέM�o;�fR�#���x��G�~��([/�"�ѭٻ�� q�}Ы�W��D*6�	$[�����%�JJyx���������A�A���d��u�`ESZ�6G�\:s��wh���Z��J�,	0���[��-�Vr'����Q�VoFU镬�<��q%I�\.�
X�9'i�Z)��A���i]�溝��5F�3t0 _M/+*@ �����Xe�w���a�e"7��]<������&���Z��1�X�=i�Cf���=�o.��t�S�K9ݺ�'76�_�BWV͉Y,t<��jal_��e���(���Bg0fP"3]@5��?������SD���Bt��6W{-TU|������m�R�D��RP%��ݚ;e����VbY��!I�#�]=�^J'����z�9#�[e�mH�fB�4�����F�m���b%Q�)w�a�=��EKQ��լ)'���W,H��~��f0O̎���[(0��ut��
(��znO�u�H)H'�̥.��Zʚ�M�⽮������)��`w�Y�
����HL�:Z_��5���v������f`ǐA��Z�~�W6����% �Ïa��U҆�U.
=N����{�~L-�k�J�W�p3�\�1U>���}�U��E�G���;�'�$�m^%�c'���i���OL�_��X�F�y��~���c����nX�q�/s�%%� i>�Y.;��ZNƂ&��I�7BH�������R4����+kY�c������,�	SK����Ա���l�����u>���E���j^J���A���k�-4�J �cȢ1j 1�-��G�w�G�M�������G9]3��.^����b��)%�<��B_�f���F5�l~j��8[���ZY��AM�&ԉ��z���"�+��p�Od����M��L���8>Z-�e��1A*�K���[�orF�^y@��h?���f�ܴ����J�HF�J�M�V��)&k�H���w���؈�+P*,#��r���#Sj:�P���׿�;p�f�Wv?_{]�(��Zc2/u?��[��N���/l ��~f���*J���jy�te��h�#��� ��4�
��w�#莩��D��f�~!sI��T�����nҋ�)��H��G̮t"Ĳ�z���~�kK���Z��+ `C�U_ Y�(���l�Ԭx�7@QV����'t��ή
�JM��C���2�)�uSP��#��=��!/7�H�����Zpo� ��H
,>��0���� O��k��}o�v:y��-A����e�8廼��	��@��͓�n
K�i��;6��J�`�BJ����ER��+�*��/@�n��&�2?� ���ktC���}�eL,�L����;Ȱ��x�ay�k1K��-Zj��ec�lT����r�}�x�i^{`�5闌����W��B���{���MT�俶����"���ȍ���]N�	iT��o���� ���M�R��T@f�~���A���*��OĤ�R�&TK[RP�X&y�@?	���o�H�*V_����0�f���+*�,*���Y-
UD���eq���M_�Ó�S��?yNS��;��S�]�̺-'es�T/qN �<�s�w���pZ8҅�ʸ�9�6ͽ�uwj��OM��A���@���_���3�������<	=^p�)V�6J�YN��0�ܻF=:ሩD�Qm<�r��K�K�6�_�7�S�<�af�7PYV��I�W���单Ўo���&�	Viz����A�$JA��E�)�.�����&����M��\��cKz���ҡ���p�R�H��:"Ȕ��L�V�V�u[$�w$�����\Q1t�rvÚ�e`�����l1��৐�L����lvSrYmTSÏ;�0SĴc*
t�~H��8�:�x9���piOƍ�����/�'$-4Jc���B���%'�fǓ�2�s���y���
(��D�Ъ����*���'g�N��H&�P�J�0�;+C)@*M�+�	�Ω}�l-^r�����Q�ձ�H�,}�?0o6�q�q�����)�A�h�J����EY[�;��Dt��"�WG�.���_v�;|�(o�0]�3�K�M��緹�Ҳ���?�.���`�L�E^ۍ"��y�r\s�LW�wι��g��L�J���?����D�A�c`NvTxꆽ��= ) ��}�䈅C�X����xI!}���.n��}ҜMFN��[ZP���|�r�gN��'����[���� ����K
>Ezԓ=���^��W�v<��BQ�_�92�R�	��m��B��;=9����ה��E�˞�i��-�D�p*")t��V�9���G7>Wݲ>-���`b�3̑	�ܧi�>wC�Lޢ���=�,��"h�Q`�]�i �]�-�
A���3���s;mPn�+	�ϥ���{2�E��;W2O��"���]�E6,��7/5�lW�RP�[�1������AofͳZ�/��"�){�x��kk��T3G��$�-ܜ��0�����)�����ި���t%���W2ܓ$���CI��:�ß�f�_��N��-P�ndl*4yb����� ���-�n�w����X���g͑�>��*BMf�e���R�2u���R���@�s��"]<YŅGJ�,�i:��vi���)����˛$�@�>��5-z���o�[Y�ţBVC��[+
��D����o�^�D�>Nl��V�c�����[B	㮕��h��}W��7i�Tu-��<g��Z�[��M����s�Z���/؝�Q����2����+-I��2`�ʠ�5`ϰ��M��u�A�&��������hi��p= 6������~�mh���x�/I�Z��º�0� 7-�s/"�j$˜�ò��]ݖ�uY*lC�d�z�)6�	�n؎�����p�x�ϔi\�����T#���P���8'����������VEe��U�Ĝ~�Ϣs��#�D�2oNlyt��g	�������L�V�$����.Hd�`� �2U�{���Ĺc5����g�����-f�٬r��@�������7���QC3#�UP����6����zG��:�\t�O�zn���y��1���>x�*@i:�ӈI����BL���I3�?�����^�\�0� ��mi�W�NKhRks��=���v
�'��'��ΙR�P&U,k��t�v�fJ��r��?��p2�
G$:H�f�LE�%�s2�^�i� i�5��bMi=bщ��s����Q�E0w��CU`vy���g�fȔ{}6���֟-��|�;���d*>Oy!{�x��ŭihԄI[Jҍ�W�N������)�����Իx���R��4���m��eNB
���#�VW��;�(�A�%��T��a��a�V���Hw���8l�=��s	t\]�A{� ��gq̀�u��G�^Z���S`G�*��Kx�A������.���.���n\:f7� ��^5&w������3Q�ل�bE���{����݄gn��>qbz�*����a��ug��6wB�Z�����[ʒY߼�����}� �(�=�z��B?S����!�l��D�qb�D���V,$sǩ��a�|<eI4vT�e����u�^6�q8W�\.�h�](1����Α�xZ�?{f�&���jc �$p�ӷ��wm��$��tTt�h�n�����=�E��\U���f?YI�jGI�?E=�_w�D*�#&�g{\�a�¹�U�>1������^��9磿Z�d�0�6%7u`��p��(T>�(BG��e��溴�d��}�����o���D
R7�U�T��t�AaL�Tz��)!���fn��]������Δ�������}��<W�t��=��x����P�k�c�A(�(u�洓sCA��餆���
oPgV�Xt^�M=�_�Bf,]��F��U�Q�N�u�o�d�oJ#�r�
[�u!����s��F����Nh����t�SnX
~�u��������V��G���T����,Gv&+N�W[�-rr�"�G�_)�S�#��_Y�G6	�~´y�i�a���y��#4$�z�Ѿ��eoiK�n����/��Ȥ\��igVƤ�N'��5�����������2~��x�xm_�y�L<�[�j9p2xlg� �˝l�U�L+��R�if�Eti^��
��-��ɚ�Y�бtF��7���׍	�#��!���&@��Q֏�ɪ��anpH��2@�ɽ�D�eF��m&�'&-mVf6�<?�yk�4���Ȅ�l��\떪V�t�/�i³��n����������h�v���×`ܿ:�Oj�8&1�4���Sq��4�*{��E�_.��~#?�;
]4����S�!� �(��l��ngf�=Jʏ����^yP��E	q{.������L���|-�^�{�E\�dK�q�c:��%Q�\F�r��!�m|�L��E�����!��#i��ͩ�֬AG���J�m{�S*pY����_r�&|ˏӿ�`��0� ~|��'~BO �4bP>z��l�a��T��%����zp�O�
42��E�
=a���I�ؤ�>�6$`3����wZ��n���
;����s(�F�E�b�C�>iN%]�}C�9=Jx��N@���-�E�v�[��i
��Y�^�G�O����d8�Qd�	���'6�y�ےn���A���]g�x!t p%��˭I�@G�H�0-�+�^H߻ܱ�%EI�X�7BOw\��X-������1'oe;�wBQ�����HkS�6��������|�L�zm��E�e_�NlR�v�YE�Qn˲�D}�kA���|c)Hy��b��3w�L�M�0}��(�E$WY:�)�2�+b�X��*I�,z3-��ѭ(s3�XH�0ŝ��h�@���ؚe s��搗�,���gK��i~A�vY�l{Ȝ�le�r�%�>3������u�Co0�(�k`����a���������m���3r	R�A7^k������e�n�Q�F�#y�[`u���C;�<�b�� ]�[��E�pXU~m��~��vt�y�4NE�x*l{꒦!�rќs�jH����9D1��:4Ӕ�f���\�!����֓�e>#���o�s�K<��È�*�Kk�Pv&[���~ϩ
�@��$yS�d��/P�9��j���f0��|l!�-��K� }nI�Vg(�15��T�Ѡ�8�\a>��@)!c�:���$�;{r����6#9��^4^�����e�V�S���	���C��y}P�e�+�M�X5�F��I�ݙ%`���ҝȠ�g&�j�M�i�����dNm�[���\gn��hБ6���)��eM��g&#��}��hb!?�S H%�b�����ȅ���0�x����ѧ8�e�#d���I�tw}� a.b��S�,�&�54����ВP��0B�QQ< �e�[�P��l]b&���ܧ\��О-H��>4!����Ay�őB����|�UϮ�;JS9=�a�Nzk�1{�Lln��",��Ս%��x�
ܕ����o�V�/�\�&�*k�����Ї+�� W_��z�UELd��ח����&�UO�n���<�ޯľ�����7�GX��z&gfН�+E�עO-�;&Z�Zq&t�	�:$>汥0�ZD4��B�!K]�V�h.��kXk�����p��e��3V����p1�\��1oξ	ͳ�]�~:�����W(�dM\bmk�������02��[��o�̞~TA�+�\L��4r�i"!_&^3��"��[BCz�L�"r'A�"}���F[I4e(�=
������l�!���Q��P��{�^�Ɋi��(�s���i�,�� �=��cʾCӘ���#����Xsvl�ɂ������,6>�0��Мz�EK(a0s<�h8E)�S���[amݣ}�\\Y�����ǋ��'O\đ��a��?&*���_K8��+�v����G���$K�FM��v��glG��Ю��,��H���`EX�	��UY�J��c~��t{S�u��rz�0a v�&��������'xH���K��{Y��M���(��x���.瀊n.�?�i9�������\mK��s�Ո�
�m�UDB���(-�f��7�J&~�d
��|�˄���q�n�N^�:܅I?N��_�(���h%T~��1�����������P��?]�W�fDnhZ �"�9�Z��m <��B#Rנk78Sgܴ��:i�q�ڊ5%�}�:�8w�[X@g�X6�|���t��$Ī��
�O P�*g�ӯĖʦr��.UE���g/釛@�2&��:%F	N�>:�5_
k�c�f�q�xf\o�����ܾ�sk�D��K&O�曯�lw(M���F�E푽<V�@R��/�O��h*9##�kM�\���	Y{�� @`�M�M���b@�j;)\�T+�睊г �P�k���Xg�o:���84Wj<0`XŹ'�:��妋� �>祂s���iB�`4��)�o/�#4����N������cv��O�Ñ�+�Lq\H}`�)��f�C��yJc�$�!,�	���]Q�6�q��� a���Z�:��J��,�J,��va�= y��8c�K�[rq�}&�J~�����T�}8+|������T
E�*��5c�����~Nw��K��o]S�4�A8����q�7���PZ��~�B�~UlO���ۥxL#�w�s#\���AN��'[��
�b���x?�@�]�SZx�`�p�Ϣ��|ڜ�qSW���w���-:,�hԻxuw���,���X��.��{J&�7��$�٨K�P���� ���YP�Bv�]��Ό���]Z�sV
h/�nl[�ij��S�u}x���2�D,������a*e��'TuY�x}Z��	�"�"�by�&���[`y�h��2=H81��Bi��X% /�qD\��P2P��PJ��D%4�X-@��(WgD<Z�(��\pI����d��Y�~
��}��v4����!t��9���h�s�ۙ��Fr�v�рӊ����U�ެ���@����s3(k"�x�<����0�F���YX�s�S�	̛Oe�c��.ĭ}����n��t�T��4��PA�N7Z��T-�ٳ�t�|�|?���i��
�!Wv�c�|�Ux�'X�
��W�T~�q��O������L�	�xx{��!���X��i6\�0[ovc\��Z~az�= �0��+�>tW����D(鄘*Ҫao�M_j�_�{�}�
����H�����M��O�h5��O�4�0������{����9n3�B�
u2�n�L;�me����v���H�fGb1T���c�O(/�����~����ȼIˀ�	�!�,���*	�m-i�$�-�?Gq�[V�Np�<I����;�w�hL� ���4��G��
X?�<�������Q��B�'}&y��/d�hN:RQ�0�cxI�<���4tQJ'~����-:ފ��V��z*'4qfA$�nue7P9�s�tq;���򶽰�Tw�c�A�@�ˑyH��r������o�kq"+��jE��/vV(�""���qm���P ��@JӴ�w��9@���3���`=c[�[O�Q���������f"o|5���:��c�S�`¡W2H�!�C$����DQ9���f��e��)9s��K9r� ЁxL�
K;m�v$������/^�6w�K۝���Ċ祝!d�qm�k��N�$h�
�P��]�<�=����[D`��62���h3��X��4S��,�'��6Y8�1�9��r��>m��)˺.�XA���:r"l'��L+�"�����1Ƕu���X��_��Z$S�����a�T�D^%����%}9�#�����#�Ղ4::��/@Ko�M	�"��1��EnP�BQѼ�m��@
�C�89̈́W�(,3�ZRd�p�^�[��ᐂ���%$u�����A:������42��֯��a��6�m]r��
�q�܋�a�.�i̬qӽ ��Y���Y�;����e��m:�9Y;�PcK6�e�݁(}��B���U�P��/ҾG�q���+ߖ��5������1"�����A������I=����9�FA0"d�r��^�Zc{z"�����>é�UQ��g�����Z�r�ł W��\ة��Vm��|�?�n����B�}c[6]�#�X�b�6�3���[��6���ɉ�=W.b��Ok�/2�NTE�G�5%]�޷�3����L���Z�ӈ�Ukd� ^�@@�Ks=�Q�q0�����h�e��s��}�CƠq��8gd��"Jf��E
:�vJ���`z]ԥ�@�>|�m1��Q;J�o�(	ug]n�l���������x�=}p��jnY�"I�.i�U6�!��=�%d�k��v����o��3*"��\�X2Q�&tk[��/��6ƅ�B�;fAe�xF�.DrJ@&���mku�(��<U�:n�� ~��W�y�∉�؁�gm0�R;Vs-�[j��u��Erߐ��d�|�zI��(_�n��kD��c���|�(��������f�������!��ϭV��g��V�̂8��c�eH���M�q��Ա��$1���Fx� Y�.�z����$�'�[4j��D�nz�������Ч��t��"?՞���B{[�I�A�\[AB��ߛ{]8u�2�������0��%������o����5�m�m���B�0�h�>[u��E���@0F�#�E�`/b��m�T?��J�v��Z����4	/��#�`�(��[�kܩ����������t�0�_��$M5��%�]I�H�1D7���؋ʩ�\��A�K�����}QL���܀��V?v,�i��(���]G�q�����A�LD�2�x󎕃������v�h��)k�C��i�0�rh�d0_A1Z��K[��W*w�Eewt���̤7�F���4���-���LTP���Q�TW�!���΄r�ǵw�F���
���PqmWP51Ӄ^���٠%��?ɟRW/{���RO�vGO���'a�=��E�W�k{��)X�_  �g�����e���2FO��_�pG׽�;+-�E� g����)�:j�&��`l�LEtg6Y!y�l�zϑ���4��M?�"����[����5_�H���8�)�]8���	�.��i�_L8���?s��V5eKS��.vfTzW�0��]Ćҿ=�9T>�;����#�^ �rnqom��y�@�
�	���nઌ1�%�j���9����Nʆ^F<݉D��/>�ZT:L���IY	��j�%lP�j��bA��*!�Ahpw�lAy52���]� B]�\�C���XK�+�ȃ���1@o 4�v��)�dc�X�#��6;��	j�b)���<�A0��nwo�~�
�$<*;��A�hCui��o����c��?P���/1^gAݭ��xlsj������z�f��~�#vƏ؁��;��@c`ᆷ���P�`U]矟݆$��|���b�tUH��7I������T�6JK�����v$^��
�<ߊh��y�����5��Pux�
;ډ�A�?��~9���,�=�Y��9� lҠ3� N������G/�#�]��{_�/�z\�Q��\S�d�g@bS�Xj6��Ӳ��r��Q�~wv�EL~�| 0�q�B[��F���R�M~�e�j�PX��U���TXNʖ�AhKI����{�[�̑ᤎNM񩂯�v+���!����v�T�m��bd�>�v|���v���G�?]o��=-֪0�xdHF�����3�~j ^��DF��`(_�2�P9��gHr���`��Z��J�3��4�6s����-�>�&|�ĸe}�-��o�!Bem�ܧf��6��/Ϟ)m��&���3aQ��9E6T�Ʒӈ���Q*i�	�?�wj9Sv��yj�Aԭ��R�`.����
ݫ�k�Ȉ���e��R�MB���g�=L�H�1�C�&4o�����=����vz� &�"2T<0�r�NQz�b���57S�����s�GD�Ȝ��!��"�ȣ�)�%���Mc�
U&�S �Μ���倱�k���Tɨ�$��)b�1T�?~{��b!]=eN4�#g�58��h���v#�qן,u!�z���Rsg��F��5Y�A���C�}
���8�H�`w`�c$Nlo��5� �C:����p��x:�?�EsB�2��v����{�C�!���m7�e�p���	a/3Z>I"�r�b+���M,�����O��bk�U.k��]Vy��ؐN�T���l�� ڞ8�[y6Bo����k=���T�[9�f�׸%=�p[����®	���#�'�כ�F<��X�{������-�oݲPv�����,���;���T��J����V��[�Uض�����e���=yq�/"����D"_å����+/���)�Lu�;�a�jvJ�{F��L]�ץ�~Po���3l+��#���
`;5����������g�X����p��nH��Wp� �A���{rk̊���`��	�<J@nP�[T��Z��&r�t�%�ʈOP���s����
.|�ҹ�l���e7����	)�ޡ��
��Z��#�;�"��B�v��C�H�j6���_�)%4�{��
��Vh�g]�:��?r;o��7�U��|K�&?�&t��X�X�c!�Y�1`j8���<1=�$b�o5zG�;{��ddK�J8��������̾e�GJ�@��\�2�:��m�-i����׫��j��Յ�F!��ݧ�,�y��c�oRDs����|j�[����_`u���c�Z�� ���SB/�ۖ�Fb��Y�lT�r�f�1��"��ǹ�O�����֘��[�Nypu�g��W���F�ٓB�ѱL���\t���/�Vf %F��n\��������y?�s��"(1DP��SW6�㟒|A��c̪m�sD����~<_@��n^m�Hz���\�~�{|]�h;�s.*� ���;�yzf�w��0{3�Ps�o0�pd �1��{�&[=�%�8����I���?�����q�
��K$���������l��t��A��@���I�[Yq%�ϔ�g��ߘ����
�X�d�mW5�l4-�Þ��`���dS����a�j�L>k׺f��[���:���!��w�^lH��L~�ͣ�,LeqiAu�-����.:�-ŭa�y�B�3���`CU���k��D�	Ҍ��0��n)�#3K
�XZڣ�o�\���,�$��e�k&P�E�D���gB��ߐ�<��1!Cq
"|N�U���Gٝq��R����l0g�?	,���E�7S�,R��n���R�����NZ6��+�Dĩ����೒L��+�i?/Ǘ�Q��B���L]ɚ��e(���Io�N��AQ��� >�? Q9��p��E� ���`���Ϻ'��	�ç�����Z�:RҒTR1�Kk�� =9���j�$=K�@bT7��bٌ_s5�MA��XA|�13�G�b��Eg<�t)�Gf�`%	jzT2>D�Q ��or�� ���u����|�q"����Inb�s�͎[�y��@���(L����"-�Ѭ��L=~j���o�\sm�f��I��Z+���f��:s�^ċl�?_k)�B�LG����q���K�Pj��lY�e`J+s���T*�!�!oHx�q���@IЧr��:�]�g��sU�Z�	�
p�f�z�M[;=��S%�xS�)�3�F����Ou�LE�	����xzp��>�eZ5`�D�������j���[���d�_ϧxt�*lm���"���P:Eгo�;� $X^,��j"�~���|��J�G���A0K���_Q����[,��pN�{� 0��"��ׄţb��&4mYaiǆj?OoP���J�Fh��ک�>��Ky��pO(�KxC�mX�j�XÑ,��m�b��S��F���b\�z������@�����=1������{}*�Cw�%��=4�~W�e�~�n���eŐ��`�*���)W��'M�W�P�=�_��%�a��4��h��2|^�������Dͪ�1?����0�97�(��"����dn^���MtU��l��������q�U����QVZ�mC�@�Y̋�����z�u���jn�St�i��rKR����I���rK�%�	uѴ�W�TJ���d)�Ӵ p?{��&	�z:��
�e���I�hq�e����ʼ=��&��Pѻ��xc	"4�d�M�������l^�W3��t���9��Ic��ʔ�K�#M5�=�t��֕�y���a��:T�FcY�J�j����Y��§Ez��k""�O �E����=L��N{��m�:=���[l��I����Sc��_>Q��+�����5��������y��ް��F���VpIR/&d?�]�M���4��n�/P���	P�O)���4���z�]=�33UC�	��LP�M�W���I�P��v��o�is�]q�F�k�-�E�2�]�h:B��^���װ�\�U�Y�&�V����i��Ø���s��F����R�,�ſ0yH�YY|�2
��s4OZ/乷D��K����~�v��s&t����U�3l'V��R��o��O��{Iڭs�����=��rF���鶱�܁D3���言�d�,���$B�q��ǀe�yL��@��N.��N�y�J�k�۾8�M��#e���!��{��#U��c����]5z��&�,d��Y�3z�	q�yD��(ϣ]�1l8����DN�1��*<��O9��:B�U�9�/O� ĸ�8���(�ꗨ�j�[����R���E�������V������*�w��-�3��G�㉑�k|��n����̫S�x��������?x���O�b�Lj�c�~��� ep9C��J�M�W#�Z��W��b�f��3ۡ5]�W��
�O(�X���@v��RH
g���.j�W�)�m~�sx_&#��hH�H"�?fI�X�>\��۾�����?g�|��){'���O�f�J5�Kl�%6�O�dd<�$Zi�fǨ��GF�3��茁8�ߌ��8�#�,�C�ġ��p�x>U)ax�@�<=��0y�/X�͂���� �q��U���Z�ΘTי�~�(�O�0���E�Yo	^>㨒Jk��L�:�V��*  <��:sV7F���]j�F0nxF�lq���[�n��zcQt�8�PP���f�����o:>o��UX��.e��|����z+�*,��T0�"č:��+�?�ɭoGnmk��G���u�nP�,Y⪞v�5���W­����W�izE}��� J��]�#�i��p��T *�TP#��%�)[xS�Ԑ�/uU�&�f,�VXc������Fj��r������aR�.�Z�;E���E3̾u�8
�#SAG�(��{�߉�j�;s�hzx B>1�]�9)�$x�%Pc��2WIʵg�i�ȇS͈�[O�年�
�7u� ���=���t��9����1���z:	��>�E���]3�?P_��R��"�]]��� c����`���}��ѩ�^���VA��N�0�8��dA�d�@�塁y���B��s��������Y;�}��Q'j��K
E`{�5���ȑ�=��JLX-٠C�b��e��j�'�qKc@�k�n#[ML���Ԙ=�����8@�:M����m����[�ӘqH`i�W�6]��M��by>D:��`�Z���CUQ�9�f^�ƴ�О�8w�[8�'�7�� {ıe\8F�]�s:�q����m�Z���|L�X�cuN��B]�n��eF�xSmE%ja��nm�#�^5�TH%q^{�X]���Rm��Z'u�y�^fNґ��1?���ϚC�󿷓���7[E��7�vx%0�įVU>�`=�(s;��6,\Z<�F9��G��Q�:�2����.�4�v�����{F��ü�H�s���`*��`��۸\b	�x"�_�1��Ǔ�Y��ʋt�1�O&76� �̯�5pp�����+�4�{D��ח)��gaTLY���l��#ُ`�U����vm�O��$�zTQHF( ��H���Mu��mc?�+" \ֺX�j��>dΉ���v|4h��>j�ɼ]��X1�6�����,~��ޘw�S�` J?��r�}�nk���C��X�&9{�sy��M���o�g}������p�0� �-���l�֜�����n���<�n��#lIs�3�?9��xl 箪D��2&�
��`(V�99�l�3�~�����lU��j?_G�Ŵ��e{��F�pwq�k�G��E ��l�݅�IT"7��]}�+%�����ﻻ���6���8^����s��+�_�����=�K�7ʋpd��.�y���&��	#R�S�,�j�H-�h�� ����J4��٫�8� �|a������X~ۨ�t0�Å5�(�5K�Ow����c˨�!i9xI����V���;��#
#5��65�>��f\a���PLM�G�hW���Uu��OF�Ɛ��0��r�}6���e��)P�� ���p�L0fuD#vE�?�B"�h�z����P����P��ˏ�?��4�s�Z�����ٟ�ʮr�٢��6�����*%=Mx>eM�(�,�ܦNNƢ���@>��)V�f���&蒸��'_��E�L'ʵ����9��כ=��
h)��YM�Ù\��4�i%-�F2�ۇ�[-�'��D��d����)k��Pe+)����k�����R��K�v���R�daE�Iɰ�t�y'��9f���)��>mO������i]�6�
3�(�L��)O܄:b �ב�H�����|��r\g�=.K�Ҙh�@ɓ��������M
!zý��>��u�R�~;��
5'� (i�A����T�k�O�2Fk?:>�-Ǵ�ɍ%�+��8��m��i������i¤�E\������S�b6��b1!IP��F�	��F(=b��c(:�Z�}z��g���Ro	s�&��u�X\S�� �e�e�q�z�5	�53����5�Pk�(l)v��P�N�6i���f���捖%�[����r�Ptx���r3d��AwX�者a۹����L�v�=�׀��u ���0��+�|��ݪ/{q���{(K!Jk�9s|�.�Ro�����#�Wv&��p�W��W:B�9ǰ�ϖ�gww�>�!5��iu���Ļ8C�J�/X�?�U_;4�$V�<� |�rj9�<�q���*�6} 1C�C�ܫ���Q�%7G��l��Q��.'��Q�&p���Z[�|�ie�ͫ�_f����Z8���]
[�s��$J���5���/�
�H.Z:�ΛBu���4��w�Eࡊ�����s��5�Va�g��kI�^��L�����vZK��?�	��;�r��FJ=Rk�p(��ڪ�qP���v�5s���y�R�3Ek�6v:;��P���/���L���bb[���D�e���*i~�Vƴ�
=Cw��ӵ�m�i5��4$�]����.$K�&䣎X�$]����ۀ��}��Z�tͭ��gIfRTMcm�)�RI��*���g��y^�L�N޵{�R�$b��V���'�Ӽ˯��>+�S8WK��(ܦ�VèĀ��N
9��],��q�YhH(|���C4�A%�"0�=@L��B�
|w�#ŃHF	���"���#�vO�g�-S��ԭ�>�qϽ)���׌�dֵC�(�8�yl1�սF�Ӣ���bK�3,�*f��C�_�����l-���on�!��A�tK[��Z�����X�×�쓬*�C��<އ�Hu�iI����E�Q@iG��Q��UV��,��گ�_(�1"�u���~��Q�b��|����� �bI^i��Qy����s���BOs��C2+����[l�/��]8�v٭4��~��R���95���G
�V�0��U�	�� �rx��U�iB浭@[�)󁔂K�{I�[�)
k�0AO��>�B�2�Ί$o">�f�����}��M�76l�78�8;���)%b�5j*��V��#�,�t����UE��wqP�/y���x6�'��E�%r�N3���-�aޟd��4A�/��lϘк1�x���FOJ:�x���3�@e�t��D�������� �@;����S�K�=����3O������O���� �́B�v��&c��I�������5�t�|J�`��#X��qv	�8�*7�4-R���1���ǒ
H��PK&=��|�v�5#2�4����O�����;Mߏ�&��)�M�_|)h�&�`�
�^(��S=��<Kr�nk�I9��S�j��Y�@��V��W��oj�9��u3��!T�\�#b��� ������'Q�s�F����Q@Za���=��e/V�ա}���(��:�gD�e1����=�|`m�}(���x�3%�Go�b�ȩ����."�Hr�|��7������jI��'d�5���a%ҹ�J;��3��<d��eK>���sBv�,��3��C끤�h�*@R��G�RLy��2�K.��`�}�#:�[/����,{W��KT,&�M��K�����YC��3�y�]x�
/�.a!nd7Ӂ}e_<)&_�aA%��A��W/$���x�/�	-h��y�� ���Ɨ��4�K�c�R��(	�#�5w-����������O��8�b#=K1Ba$��0<m�X�E8�T��^���N�ȯ3jd��8�䉩g����*Y�R�-�#����@�98gw/��ݚ�A�&GO-�t��aqJc���lcΚ�f��@
�Ab#:���|j�DP]%���
�£�� �׃�G
Y8��������A(�p��)���b�u"7�uJ^�>��u`�(�D���v0	�ݲ� �&F���]�@B+f�����[�V�$c�]�k^'��j����{%	Q_�P�Em�Gk�d�v��h`��bmfS�Ɋ���6���U.�����<�����rq�rt����0B�,��0�F 6'	����T��P#�~��t�'i�E���%��)oЂ�J�~n���A���[ym�Z*Nn����nԁ!M��讔�|ݝ�){S)��`om_�v!IFJ�&���Ο���{[�x���'Cc��:tMtw�!TfWbu�v�'���a5�ץ7D���#�^'r�R�_fVM�G�f��we��kJY�iP�fN6eUTs�/�, ��k��޸�ހ��xa}�9y��GT�!6"�%����=6�'ȍ��]TZA[��_�ע�3��%O2B�FEBg�qej@f��
#�F7C���oM�?q`�EȮu����Hl ˛c�
�G��N@��1�O�A���WbU�����?�'��d[��#�#��͞[��R���J��D��݉d�������A�!����őx����b�,͈&��K�v�^VPF�,�#�����_��#&Gُm����}�1k�y������`��L!C�T��8&�FV 1O�ާe=.�M��S$/���j�+h&��9<
��$�F0D��S�2%��7�Ʈ�W����Y%Pt5��q���$�j�'-6f�jZ������c���O�O�p�`�:��O0�)��~�̑�G�[D�،"�w�
,��|q�L®�ߩ'l~̚���q�W��t�$���Q~����J���}��.�H�~y?���P���|���Ӎ���[FYk����,��+����-�(�@�$�0���N>�[s7/<�m�n���"�	��S)��0wTmfeyX=S*��*�!����^4�F����R��f�z<bj�5��cc�	��z�U0�������ԁ-���yH�;���:b���n�u�����*�U�����凵�n[�P�����tOt=�Z�P*[��:�KFGJ��Qtz�>�mG�_�����7�],M�-����.3Dee�}�YWEu��]P�l���΋\�%���V�ぺ5�+��E�����U�F��J)}⣗>lMe�)��o�B��s�i��ɡ�.�4OMg��̡���g�����l�ã�!h;��%�����T'��Z\@M� ��f In�䘜��uq�d��oÉ$T�U4�CF|W	(��M�ܼ��w� ��
O8��5�T�Z��xgϐ �Jg������[w����E꒘����*^���g� v�+��6�Ff����N��R[ނ0C��o� �T�Ӯn�9�6C�)�5=�P�
���ֈ@���il�E1j����"����TU'
�V�eVv����?��a�u*�@d���yR2�����J��l�m��,�s�ؿhi̖g<�����/ m�<A< �Lc��@I;�x����}H�v�����O�l��RX�Ŭ@��q�����Fr�- E~Y�wVa�`�̇���W6��,���(h��q��L^�:��Jg�Y��ȴ�t9������V�&�ݴH|<�K�ϲ+;�h�噍�y�t���#F�#<X)+�~�j?�k�`�����r����~���)�!�R;�OA�`�F�M�����j����>P������ ��/�>����	dQ��2{`���SU
8�kD�W�J��%d8�/�u.���U�Q"'m�ɳ�|y�B@O�m��Ra�i�ay�۪�9��a������'t0�0[�tt4i����F�������}�C:e�X$wa�:2�MY/S�S��u4rCgV�;�����sNn�ӭ��{}$���l1�z�3yw�3�i��;E���W?֭괅0�0��vp���a`��s�̞�2 �.�/��)�կ(Ņ��� ����`oN^3?�`����������݌=��b�<(���}�ң�#JS���9��8�TSw.�IQ��lH��k(�c�
yP4�ۘn�ְ�D��a���}?/� ��q':%�6��hD
�w����J�O�-Ӹ<���j��8K�d�A��Fǀ��Y��C��D)�j�eA�96�V�=��SG���r��{���Oz��J㐛Ho�uٸ�	Ch]9P���*��º9u��<��i�ۚ�ͻH����g�U�%6���c͹�!��w/S{:?p=]����BB��=�Cd�
Jq������9��� m[�i�,L��c�e�{_O-��"T���ɑ�����Z��ڑFJ�]�I�jR\YY�O�,�*!��q1�4G^��c���R� G����y@x�������.����Dr-˖��*�R9@�>-	r@^�6���>��n'��l�D�	,�+��Vz2�-؞���.�=�ѽ-]���s���]�(� �Q#V*�,r��
'Fh�]-�RY��i��X���_��)U�P��K�� 9�a�:-h�f}�@��Kgh虎ߡ<,�r���x�4o?����I�2Y� V�}�3��D�Q|R�/�]�$����'LfJ��[\������#n
�k�䙚Vd�i����#������d6�]JE����k�k�����V�i�y�+`3��A�e؟��d�J��LPU�Mc�VƸ�L��Vg3�j,��:�j(�] q4�l�"V��ZBۢ������.�~�4�ڽe�|Nו.���ܞBee4�npڃl���5H��	-w�>�nRg�lΐt8�p�(��+��̞c���E��ٙa�U�D.Yꞯ	�l��h0��#�Y�x��AP���Ř�Bƿ.OQQZ g����i�l�
H~U��KX�f��ѐ̚���,�㑺'M%Y��pʷ�>�ȧ0k�T�^Z��u��:]1�`h"���T+�d�ݔ�oz�Ҫ�Գ���{�+�t��	aX6e���Jyj�)��њZ�~Nv��i��2Y)��s����:,Bu\� h7�y�Im`��?�w��B�i�Ұ�7���b�O��y+��>4�ȁ-��}�p��9a�JF{��lx�9%��UQ�O�:ɕ�*lyI;z�5�:F4����Q`B���ٕ��ݤY1x4�|!o��R�B@H��<+���B���K�/a������v��s�䰽�s����N���1����5kܴ�����߱�|��.
�G?	�$�4��D����� �c�7��ə������݃u��C�S��%wh�������d0�u�S^W���(S&3����c��'����	Ǿ���4���3����t�s����'dC������w�=&(���/>�E���mE�dM��sA&�@Q����ax���0"k���1�yW��,�Ǵ����r׬��o��^ve�\2�� �2SbkW2]����W6̬}�W[ھBwl�iJ~�.Q� l;~X�S�		�!�B8�9V9=�.4`�����ά#�y t��:<k!�:�<�x��b@U&|�s`�8t���(u���//ġ��9!	+((�\��\�j�>+k�9{�1�q��	ph'oÄ��,!�p�������w��}�1���:y���0�(X���L�*�0��L���P��=Έ����܍ݱ
A��'�������k|��`�Y���P؂�fk:�tvJ�����{$�Eɸ~��@d���P�J�6��v��ӽ}�� 7��c	�h5|5ef��
zW�ԭ��1(����е���X�����d��$p�?�
�|(Nv���i���n+�O�-e��\��M� g�\�ǝ3�>uv���>�aM�:�9��E;�#7���}#���Q�y�h��ǱpD����*��2-(������GĪ #��4��<�C2#����C�y*�P<�3��*os-a���nȍn ߢ�h_C"��j�����~���k��)`�N{1�M����f�����၎�\�o�<�պ^�����T��}\<�c���E� �dV�B*DX�5��$m{ZkD#2,����	#:;��=m����������̃cdL�i{��@́Wk��S��y1��H��h�IE`I�JA�<��杵���e���OMil�䤛��
o,��������8�;�	����'_�p\�ܬd�{���]��"�\�.�++�+X��,6F��%ڔJU�O:�	`Wr,,m�
�qƶ�_d�fQ��Y�Gn�A9�Of�U.��/)eId9��콢-��X�0;F�Yyw�,����;~�޷��E{I�@7��䃋u)N�4N �F�"C�����*��T)g�Sըஅ�V��s��J7l����QK��D�B)a����p#����EP�����s���Ʋ�=��50V������P��^oЀ�rji����NT�+	�
3��.�@��	�)OrB���T�t�ŉ8��|DVm�y�(�'��3����y��͕.X�%F:	!�M�ۗL�WS�R��枳5���e��HJ`�1NC`!<�.<�c�>��4�Q̅_K�}��*��[��CB+ ��_H5�d	4�B�ɳn�ǵ%s��B�x�얿���'��o,��q��ُ�x	JD����￦�5ˀ�>�ྡs��,%z�5�����)c�������}շ6��B���
����#¡�9�dr&VR> ��F�9�p�8�r�#L©��|��0rG���)	d�i�6W��5� �_d��a})hȆ�i*�,1����f�@�R���̧�&��	ʏ����i�<f
i@�`O�on�Wb�VE�A�Ad5T�F���;	�w���Ȼ���y�Ϗ�����׍�m�|8�u6^�{������t3�e�kQv����ώ\����r�n�y�,L�/����a��	��S��M]��c�����w�1^z�Q\�9c'r���Z��)�hMB+��5sMI�5@��)	��@��AZ?-X�DG�s)!�PMNO,�����Y+͍3�n6�36Z���5��l��T����F'qf���p~�ݙե�ad�"�
O�V��+���o�ڎ\{��������6>(x�ڊd����6Ì��:�u0Gt��}<�;:�lQ�xؘv�l���F���m���M�(^a�����b�o��-|m�c�`1���b�XA�Qx����7�W:��~{{�G���$R����s,�h�����L�=��'�����1���@���{��Ņ{��ej9@�00��b2���r1`����ڝ�)�ߜ��]y����{����L��I���$*3�'�F2�@��%�Ӛ���~��f���53$�ÝymG�l���؆c|)��Eh@����1zp-*
A�$��A��0�^F��O��)y
d����{������ˮ�MG��"�&:HM����N �Kl7
5�|ȓ���NqJ�;��Ɍ�!W��~Nf�6so�dʀV��MiH`�S��3)��{��m���LcV���;92��@�(<��)C�,�'�yP���ȭ/����_3�.�Ԇ:ӽKS1#�D į�^<���>��|dFC�2t�,"O�z��k/ӝ,O�b����� u.�	]����cŁ���WF�v� A}��6�V|T��[��б�WL�i�� O6Tfq�Vt�r���)(���RvüG}b9^LO`MLg#���Q�R�c�pA�p,�I��(ke#7�l��	u-׳�a 	[;S�㞩 ;��a��8�z���p��es�+Qe���O��x�]j��%���<��0Fv@��t��rƫ_��w1�P��0T� ]�y]��\r2�̊fKJ���#�{�0��	�{v,Tv-�����z�C<�M>/��S��&��#�n���aW[R�Pa�������L���8- ��������U�#��4d1b�i�S��0�����ӭpq��L��]��Ae�tͷ?��H
q�0v$*���,��p��z�d7-�[
p��(�I\̍W�%:��Cc9�Ϗ��h&P�e�Cl�{3+U���%��
J+����A��T�ru��ü�#W6
�@��6�T87�e� Q�`M4h�?Љ$���V
W�M��`�(۹Ȝ�-\�2���V�߀<P �n�W�1��C���^R��c�d�~c����ɛ�w%��O��TCJ"�P�U�K �fWP�� ���P<��t\�;V�B��]��=5�IF(����v7�Z�+����	P�������s�>QI�;J~�0�Qi4�;���!:H��SE����G���O��#+��a�&�q&-��!MvqB#���KV���L�ό @S��3[/��Y4�A�ߣU��*��#,��A��Hj$}�8<|�t�l���3Ё8��O�2���]������{����%M���dg}�/8��h�ȉ���R�im�PI��ܳ�;"������6ہo��xAp�UؚcPxPn���Zy�yG�*���'Z�`�;�a�RL�1���;�b=�s�\���[���v���~쨞� =~ݞ�F.|G&�����ɈDrD��� �+<ѵ�Vn�ݲ�t}HНkUu��h#��w��%��W�-`d�I�p��g�F%�>�7f�s�2��Ħ���댒�q���U��ҋ�ōz?�$/FAL��߆
��J6�ۖd����uD���V���ű�^�K��"��uIr3h䧣cO����UT��U�l;�cWV���:H�Z�D���\"Ҷ!;.��w_?m��]YU������ .)�,����'�d�sD��#�l���qҺ"v��Ep���0��8����� ��(�IFO�9vٰ\�����u����8�Q�n�@�'6H�<KW�]AM��amw"ጀ3�v��)����V�3Es������v㡔�����T�w�e%~��U�9�R��V��'.T�;�)��8H����I�{��ڻ%[t�>��i�^�iL�����\�����)��TJ9�G��|�+��������1�M.���_:�|���O}��{�dH�V��k����q�^�������~�������#������Qb�Їi`�	Q9��w�TCz��LK�����<n��HF׻L�%ɇx�/����(Iһn8,J�`��g��D�`7��E��	��$�
�.�<Ͷ�:E�k6�z�.�qAO��dҝn�avfz�,�*�m�r� *0�H��W`��`
̚\.�]��u�"��?�hF�d��,�gm���l/b�&Es^��l�Ւ3��L��+���-B����Q$x��k�w�n��k�N���T�v_��a�*]��=���<j���.Q,��#�7����6{�/����� ���Gk��)�Dlu9�xy�������H���l�YE�R5�h�bb�	�_Ǽ(��5���� �GhE4�:%�d1T��T�%T`:8+�5�y�Y���v�Fό���� MsC�R�I�YJ=O��Ra���
�5A�s���7�M�VO3�o7��E#
kJޫE&�_���qw"%�g�rx�
�Ƀ��t���Q)t���5aWa��p@�O�=�捒�G���44y=Wב��^zx %�*��l��[�KOR,���u����v�%W�;cS�A��~X���DUK�@�^��bq�)QNڼ�X�t1#i~|�յ�Ml�@)�{fD��!�a��R�	E��:\�z@��M/4��n�1
���O��:�y�KVv�o|[w�@(��ߦz���������8e�&�LwS��:��ؼ��Ou�|f��!5�s>��!�?b���U��zC������ޝ��t@y�w�7���.��F�[~��7�P��⓹|���6t��	d�A���ƿҙN���Ǎ%�C���v~�*� 0� #�$.�0�@��	4I� �.���'�p��OI+/��ԭ�n�G��w���>@�5�>}n���. �ބao���!pzv����h̪%b��V�M�ҽ����A�ư0�S��䆀��-<y�L�f�m6�G�&�?@f8���c�!�NEKc�V��7s����V�u|���Uۯ�/ns�nZ ؉��y���韭�x�c�gbj[�4 E�����6S/�+
L�y�e��H�B�8�0A>�>Gc���K[��ӂ��m]��><Uf*���ٌ�+�WaX���/R�'Y;�U� ���z;H�ȹ^(�yv��z��3
���*��J)�܃ͳ;�BX�ց�<~�s,�ۆ�
�1Y���|{�|ٞ�e�ڐr+�G\� ���c-����d����?Á���'����Z"��rp�j�&?���<����o6����}ί<���C���E�ՄL��<�V3��K�:z�����(y݇R��4*_��P6t�n�#-�\琲�rea�A��S���WX�=�6��K��)���k2�k��
�♆����~"(��[�C
+���+ �=�u��fsqmZ7='[-���� �(���J�
Q��\�Mw��b��+a>_�K4�����7�`ſ)��/
A9�&��kFu9�8�� 3`ʮC𑺟��)Nx{|�%�̗�~�u,�^q+}&�ϔ���S�ia(�.>��mH}����{�rA˝ň�ß��fd����U�xz|0����7Z˙,�ww+g�@�g(�U��s �f�7	Q�T��5 ��^p���$N"�4�����Tf�}5��u��`0=ߝx.��y�������zw���^���#� �+{�Z���rE�@j{X�^#�����ߕ[*�lplT��D�ζ��fBE �##�Ya�X#QiǓ�Sp��+#���
˹k$��Pv'�����9����_aQ`r���qSn��0We�n22�S��E�ch�&\P.QmSA��1�F�V�(.���*� ��oUvƐQu��ױ#/U@G��HU�Ga�k�=V�a���ʘ}��Q�z@���c��d�%7�c\W���4��o�C�b����
���`�f%f��;^"�]�)~�5��F9X�/?2�ݴ�c��9�ΐw���ce�6���5��鎥'��iu�;4}������*})+R��?���	���Ξ��h"P��On�
��dk]�9/�Ln�P�\q�𸴇[���	�P>�eY����Ѕ+��h{�4�e��4O3�:���AX@���)7��V��#�,!Y���4N-¯������B�P��e}Ο/?m��:�'[j�,E�˒Ό�. �.����Z��a�v���y�[�q"�1v�� g�'�n���r��:��W�ȍ4��r��;�a�hw��A�b?A��.%��2l�EA~V���o�P��꘠��j�L9�F�Q���KKu��H0Jb�-�(�6~�f2`���%EW��k$v���N��������ʮ�<�R��Rf҃�NN��\�qM(�h���4mƯW������)h��40'��t�l�*:j��0H=����	�� j��x��Y��?��{K绐�6��T7r�r�]y���}�o^B� �~��ŰZ�%�ŝ���@a�L��.�jع�7p����ɬ�����r��bD��mC)t���vO��(}�[����!�#�U�`|���.3d�9��r����4~Ey��+��ʥu�?cǮ��G�� (�4,����?����?{n����ӡz���E��i�\6P]N\t�J�d����tz�_]�fSc�X��K��<�;8�˯�Ә`'���t�U8"�#i&8�35���)b]W�!�8̗���-a��;�&��B�`h�: a������E�){ӹX)Z�%�o(���S���Δ�a$Չ���0����5��9�H%KMq
Ϙ���7��W�?[�-}���q������ �:E�:~و<�����t,I��ɏU}J�����h��g;����V<������zd���ƀ�:Cʠ�y}wg�'���dD�8E}ˠ��z��z�B�W��F��
l������b��	%�e@�,�Xr5���R��R�:�՚������-���H>D����=����&�
�|�F�BB�r/���d�x��.$�S����,Q9�4���<Y+ץ��K���������o^0��0��0�%�M`�p�Mǖ�[nc����r���ǫE�I��wW)��P)�a��F��tS"|� �����E/�J����3y�.l����=(���ώL�|b�����N�gR�����ʵU'�{/�����]�6Ąs�@'@�PXG� ��+X1a���2���4�ώ~�B%UXx����vp��M���	���a�q6�G��R�~?��&��ܲb0�7���A�h�=�N�d����%j�xΤu>���x*���z�E����#�H�O s���Dt&j�e�x6��
V�foZ5Qx<�=g$��㲻~~0m ��D٭�e(0�����}��l���}smW��庘{Ф��N��j#�'��bl�'% ��*S�V��IR��+�~H���"�ҫ��͑��*��� v��>����\z���� �7���TH��_[A�z?c�4!��ɠ��5ҍ�=��_�}��������U_����}���1Y:Cc����,4�ki�?�2�H9�>o��!OD[*�a���ק���m��L(L#`ze�x�l��a .�/j[f�Yr�ڗ��[E;�?����;F=�ו	ᐮ��G%��+~wz��Q��Έdo�n2�x��fS�a>:����!(J��%K�w	���̟��<N�`Ǎ^r����e��y�C��7��\�^�Zc�Z$M��k����q�6w���u��m�W��CѴ#�P}	Jg3Nm�Q�~��g�qT#�$Xa��3|~�f���ͺ�Kt�@�Qz*�����Bm�L���|�.MՒ�gJ�kם4�A;�m��7���TjlF�)��y�^H��q�M�\Bi7޶7/�JxO�wY%��z���n�մ�V�<JG��r�hA�F�=�����z��7���7�ء`�(	��촶Ҩ�Q�'�]�'|�w	5䅭���rfw��-��m��/�i��z���M��j���D�e0�I4��oI�ؚO���Ծ�JD��T�
F��E�	]r�2$#F�_�"t�y�ٜ�8����:n`�j;a5��ԱVA&LzƔ��3�����]�G
*�0"��K�����ӆ������J\@�P�pXc��Y��@_o&z%�y�sw#Ew��?S���н�-�1�iE RAĚ����I|-�0#X����?VX�-
Y;7��/����˩�[��q �O#�B*vP�A=A��"�����vw-�u$<D�ur�C����_�[�����C��D�_�)�RM�@���7r�\�&�e�Yqļ��FH��$�ցmw<��C��O�e�2��M���>9R�5�W:ZQ]�;��Q���G*��{8�F�ʢ��y�/�l��)	#1��3ξ���j+'zR
� ����9�m��_w��Ǌ*N24#\�y����&�q{?HY����Ib���f�pc�=���P�u H�b>N����M�Kr�><\�K��^�%�3����4����� 2Pm/�!��7�p.7��|��d�o j
����"p����Ƈ�d�I�Jz'��G&������Us���z��s�EM�#�0�e��]��ctC�W'��J�e��[�ΟJ�Ԯ ��ʢ�sYJXq�]iK0��&������Ms�9/�۾#-A�Q��Z4���f\�B���ɛ��U��y�����6QRݾd�I	��G�kS���7��v�Dư�'�e'��y�a�����'�2o$�&�#Zb @d�����9����?$��p�#r�&*�p��Ѓ�[&��Jget]�P7�5��_���ۅ^y�N�X��Uh�c������Q��Q���Y.G£ fj蘌K���s�VX�-E�E�N���	�@D����bqqh�ƌ[����5ܥ�~����������'��~��zM$��
�0 ����f1LN>��5��e{p�tm�F��/�I,S=�L�5G��=."���Woƙ[�P�^t?�!I����&�����-�j��s����E�gM��D��7��n)�
�Q���+p"��Ak����}2l��=�s�bz�pdB�9�^f�^�>�8�ā���lz����s����6+�OA��=��Mb+{�s$�I��X���B���;5V^&\y�	����ƿ�Ths��=���H�IZsܒ�!���
%�0��Z��+$j�䪙-v�w\��ə�)?��d���p�4[���a���|ƞ���Ȧ�g%#�juY��G?y����]���KX�[M�?�};8)�P[z��iiEX�x3�F�}7 ����yd�898�+s�YJ����I�C\�G<�PO�����>��m�c��M�ZX��'�o�����Mu`��
��Lmx���%xM�ە�����Z��>�6�='Pw�c�Q����x��2+;����jȿ�3�V3�Q�M�י��b�7�e4*���m�XI�kJY4�3��}���fn��f��f����U���~+AΖ�̂aS]������\#`Q>���.G�JtU��g���J�Q�Nt��2+:3䣌wv�J΂�؟C�.�Â�&�Ϻo�<�K���c���8�ab�c�1�N�U�J�(^!�Q��D�xn��Yw,���cܔ������ ܑ��&�铊t>�O�`�f�qa!�z�
�X��"�{i���CZ6T@��b>��?lU��%��+���j�V�=}9L���JR�.v�s0�R�z����̦�ý��EP���?���� �8�I�hν8�҇J��c�9gK�E�XE�(���u;_����6ɾ>�^��ev�%X��x*����
��6���k_�V��9�cb+O�vvw���"gO�	����Qrl���Kŕ�)X�k�y�D��Nk��sBA���oYT�ơ�)�\q�}���źrϻ���b�l	����Ͻm�3��_��M�5�|�{�+/�:�H ]�M֐/?�r���<�d���Ӊr)|���u�@����H���*WPk�`g�C�\h;.bo��"�qK�5�?�C���?�4@��p_��	}:�dJ��ne�䊙t�԰��:�?�75��Z��Kojw�2q���Y���E@(���Uq���������k�lG�s�E������#,zڔ��j�������Fə'&B��L�C؎��VT�0�3'�6e ǐ���[�L^�vU�
�aUH	UKy���Q���/�K��^F�-׆|�y#����9��$	cv�O*��������J@v.�A%����<\ޠ�E�P(�]��<r�^񰏫p<@��sk��Hڰ�F���ݨ�6��]"Y�Bl�T�},���ٴ�.�&��L FL���튝:���},sFR��4wR_$�gz>��M�y���0��e�ͣ%Y�(^79��*q�|&�aI��{�||��i!|!e�����;"�����t���
�&sB[��E��I�(���䧘)P>���h�6�q_��(��Ǩ��h�+����x�FpE��F�F*�lq&)Jlr�D�n�,��������gO����Զl��?쓏`t� �١b��j}�Z��g[I܈{����LcǾW�:��c���̤���G	~-�u*5g��Cy(`��O��e���_6.��ŏ�M
Pt�I������S��v��#��;eo������<f�C�9�4��Hw��O�4d�t�ɦu�����K�1����������&�G�����
��V�ޏk"�xE�K���(�B�3����x;/z��u!�X���o�ꡇ[vWf��!N�]�sڜ��n�d5�Ż`㮞FF�����ʡ=_ +��y/o�Q�e��F��L�1$NS�6��k3�io��P�����i>����cM��۩��4ߥ�j���;!�Ʊ�W('���|X��H
��8�� {���h���C��)�3��hO��Hue�O���􏽲*�4f�g�ԡ����y�ϒ�
��˚����+���%a@f]=�:�b��0?&��HT�$q�cJ���2t���|4���,-���"�B6���2$�����d1$H���䞪#���������S���c A慶C����|q�k�t.���@�8��Y���]l;�=�4R�0]M&�*0l��Mc�<�U�!�t�Mm�]��(�k��:O2�m���$��Z��N��a���q�6�^������^�v|[ɷ?��t=����r�ES܇?�T��h�&0��;�2���:����u�Y� �d�i*�1��qr�$|�V�.���������X�Cʺ��$92Cvr4a�?�ª���8�^����岐-��0�^H��e}t�����Y�>��|�
ǮÕH�S��"G��j%�p��;� ��oir�t�����N>W�	�F��e(�ǣ7dB��bB�Vi�\��ҴA�ٯ��6��� �ޞ���[xf�RI8�FEoDo������"�e|�}m�z<<���0h���a�~p{;��r֧/�O�ߔ���b�cOb5�
���f��J����@���ʵJ����g�s
|��4�M����F��(�)#��'�0��Ж�kk4�����%œly��"����������{�xq�T�a�6Y�22���{/!L�c����}�Fy�ܞ����\П�ưǧTBL�˪�7r˫<�'��nCMk�Io��.9˜)��ӿ:q�1N�(��ԧ�s����͒�G7�ަ���|��Y2��Y�����"ҽ����-����[�Y�Zo�4}�ύ(���"͸93ObE�z_M�w�`X9��m�� �Ϫ�2-�o[9^HN7X���,�W��g��J�x
��:t��y�l�W`�'�hT_˾���ܪ��I��bb�"�aR�s�	Bj߽����ɠE��o����ѽ���B]puG��%�fўVnB��9���J �{B����-<خa[�{ +%[_���TG�Z�*4���k�b`K܏1���!F�����3�~3��I��r�C�\<�8��T��V�<�
O�x_pr͟%9�G�7�-�D�E8��Қ�b^ܸ��(�[&L����Yk�l� ��2�"|}��,n	�{�o�����F>`��������K��U�Yk7��h>;ĆA�-��R��(�[�#j"Ej��6<��B
�[�<���r
�D]xN��p<oۇ߇��&9��q��T>�w!(�Bɲ<�ewC,G2�A?2�O0e��L�8T�걮6�J��l�r�l�~�ג��Ф���}DJC�R�e�82~8ژw�=���ʑ�fvy�*��6����j��9���xA�D���YO:.�[ۦ���N�g{�{SE�v�����Y�d��ӄ���E�	���	�r
�����O�RIk�]����Ҧ�'��z�\Y�N�d58�,ѯ	�������6��ߏ�ݹ��~ҞG���`}�,~]蘔+���WV�j�r�~2���g�t=�WE C>b��R'j���*v��$皧�%9m	���9y�>��A����<�����j��m(��U��,{9>�G�b^�;� �^��1躋鼓\�����y���JqVQ�ԯ�>tq�����>�'�7L/U� �9S�|�I�`j{�3�I���eԠ�;#45CYE��ߊ�����r!��䣨$a�n�+mP�����B�l�c0n��'8i���s`��.�"TſS��zY"�ЉS@��]�ab[l̟W��[k�,G��J�=-�=t���&�͖�=dZ��2p�kI��w�%њ�T���Ђ�AW'�v5�Օ�ɀFZ
�qϭ|2����"�6�8�%�wߗ݊0��� ]����%�� �0�.ܐ��	��� h�� �e
�ut}`�R�'��h�~+�������zѨT�ڤw�"7ӧ���ԣQ`o�?�Q;@(#1sr�ī<�>�$�� �K�,�& z�"s��mF�q�)4��4���!�0%x^���b�ح�d]�����60+�.,{�܏#�����̫����Y�c8�5�����K!��sL��D�^�6=����!V
O�E�_��k�[��]�oW����2�c�RB1�#�5t���a����Wp8�os��xW�0n����SF�, VK�CU�o�Dt��.���$�>���SM
3t�H�s�i���
'W���� �;�y$�hx�Qn�Ks���oV<��ғ�\W})��,�,�#X�;�9��eC��^pr��a�t�Skq6/���(|/AP�Ղ�|���Tj__9	�"އ������4��h� 
�<�m�� D�M�-�|��\C}��<�~�����R[�3ë�a���a"F���Q΋8˴�A3v�p����!�GՊ*0�t��0	!&�G����~����}Kg�~��DVD1cP��7_!v�U�S�$ʘ���`��K0�Y�g{�%?���z ��9�������sئI1�H�4}y�,��}���ӑ"�O{|>IǗ�.O'&�,rmHӇ�R`Z+]*��z�uP�xY��'��?&�/��f��>�)�����k��3�!�xʮ��438eJwڲ��z9��4���]�p����qed��7��%.W[�S2+�'v��ٶ��X��RG�r�L��-�)�1���շ�<��6����/�;e]C!��5 ��QG|D�63�&��Zf0�����K��&d1�cđ��wM���uo�V������kI
X�L*_��ظ(�G�� ��:�C���:R�v����7�:��e�#Pߋ�K����.��Y�-|-h�{�,��[(n��-z.�{*�952�#���ؗ��VGt9�����,�k�X$'���6�B�9��'zoI�ka�;�i���'��T���Fg�n��٪[���-���L������F3�Q�:�D�T(�Fby�����η4�3-Ɂ��î�����k��-��YG$����C4.�xጻe��;�_7~SaQ{@M��)�O)������.r�?�T}vi8,��D���ن�qb��
v�oÃ����8z�\1�"j�QIF��(�̴�N)�-=�L1����$5L\KLK �9�*�k�Z��)f���]�z��Z=���.3��1���_#$���N��@c(�q�I� �Zg|���L�Ԯ.9����L�$���P,c#�DV��{;RY`x�G��I&�F1�g�⾴u��wA�z�k�`4`ea�}��*���BD�U�Z�W4W�s���F��I$�g�3�l��T�Úǒ�ta���G�R�=���_��k0�i�Y����.e����[�~!���3<(��/��$�i��g��r2j������ �L �t���~��w���=]�Lɜ�Wg��=� �w���rfʪ�o��;6�8��J��&�7�>%�U
�`?����~���`��]�h�R,#�`���ۇ̩w��1$�?%;������TnW�a4IG�b��u*�]	l����k��g}���FM�rne#Ad�1�^�U\��zX��D��M��v�G˖��l�y��bD����r��o��RΫ0n�����Q�֏�j��q�b����7ϞB����#g�2զ��2k��
'�����6��y'�8<�Ԋ�h�<�/����ݠŕ���h�Y�> ����d��&#�	@/mє�h&� �~�p�̔E�R����~�wm�d��?�[T}TO��u�J+K2Z���F��3����°�M�8F�QP����՞���0��^z��f�ʘ�LIq�"��.rm��8�]B���&����B�Jb��·��Ih)����[f[ֽ�[���É��_�c�&0��ʁ.eu�<)+{jƠ���G bޚ�wbk�ʕ�{�yXJ����>���%¶i^*tg"�)Α݌��ǲg�g�،z���_���Ro�^
Y���B��<�P&��V���� R�\�)-0�;����j�6��=-����VH�N�̀q%n��`]�{���h��񜎝�<�� X/$�Rp��F �Z� w�at1�P�	�5S)�z���%QWD+�@�x�[쮏&F���qj�B��[R �Du�6L�^�1�pϛZZ!�}��Z�\�2�?𱢇1���z�����}u�\���ĸ�ظ�q��޴5�R'iJ�&�C ���Pň�wWW)|K��B�Ѿ�I)t��TZ:�m7��D�c���c�q�^ʕ�`q9vc�i<�#����5ˢ�
���Y=��<'�Z%s0y��ƌ�%��(Sh�o\r
�?WWѸa��Sx�n]z�(n��.d�f���\�NpHw�����֠w��M�r~�f��lV�"� ]n���T^#����%|$��'�W�F���j{">��g��pd���O%�q���)<�t���_X���l�-���Q0(���$iI���W�Z&�D U�Y�Gw�D!�/&{ot)�ֳ��䓫���P/�)�X��װ�F�8Z�eh/�ϟ5���$1��X�8Y�lh��Ug��.5��]��u���̺a��
%�P�	�~ �v�hF�~y���ᩛ2"��%P�jk�Ǌ31��`2}����e� Y���VO���y� ��ټ���sP�w�VG��RikYA���	����P
�K*��m8Cuw��[���B����(�{��o���9��6���*]��O�E�N�0�B���u����y��6䇒�O��폣���8n_3Ҩ��x;mJ)��2�X�8�C��$13Q�����G�L�ǆ#9a�X.ߡ*���
ٯZGЗ�SN���Ҹ ���z�V�y�Rgg��o!'��b�H���d�o���j�^��ÃӇ��: ���t�������U��p�
��%)QaEc�2��i��դ�u�#n��#_��`�ӨM83�ņ�C�Mʝ*����Hç�9��R:%	[�ԯ�dv=		.��/A��`�],b��}��z�Ѧg�S4^iJp>���Ca4 �q˪*��G��e.�z��W�"���B$g �R����Di\8_�p�M{L-������P@���,�~�V�!���=��E��!�᩵��H�����ơ7+��\m%�dc�s`x���1JyN��L�#3ؾ�- ��4��M�7'u8��RV�E$��7��H���?��������}ۦh� ��䴋�|�Z@9�B��etBڠ#*{���d�'�D!Tm�۹L��J ���-�)���#���6 �N	��d"��e�I��҈��!:F��;L
���Æ��u�n�lN��I��J������m�Kꂩ/w���JQ���H�Y+�nO^i�"�r��o��ο*&ι8�ъ����t��US�-v�`S���^�1h�e9�p ���0E�%�[n�-�N�p����H̑
�c%���@q���J�=�1�S�+�a{iPO�ƚ  O�H��KQ��ᘂ�y̺�l�?�>%�K�-;UG1�k��`�y,V�
����F%g\Q$�Pݗ�=?@�WXe��B�"�@�g�����س�-nHY`������)�CV�\O�S�aX�dm@<�a.���������n��觡� t툰��?a���A���Q��I�-y|���M��-�&�l�+�i��_�v���C<q�U�6c�ʜ���Έ
KŒ���^�(�G�v��$}ʳؠ>��zU�����]����B$�
����z�Ջ��o}iHD�3_��hX�{Ml�xx�z��K22��ƝY�Y���C���v%jGP�daH����>�m{y$3��KƷ��J.8��=Kh��i>?�Ȇ�;�����%�;el�]�a�{�����#_5g��	&*Ad!y|.�����Rk$�2L�L4W4��[4Ao���7��N�ί� �2��E\4\�4����"�6��娨��c	���=W�j����Xr�����1�_w_��1<����}cKs#�_�q�Ѥ�&�5t@���q�ku����b�2�w�2Y��*��NQ'l���������yK_�v?��e����\؁5�#�f�7�>/C���X�S��dƣ+�+��̩R�M�&D�����Ūã���.ڟ�[(y��
0���P���л=W糲8�c(�� ��J^�M�ӥ&�C���mX��_�7��uX!�{B����H�u�V��ߴ��]�z�L��E��Xp�|����6i g���2��:9ԕ���eI��'UWq����d�엝3��Z�
�	d[Q<a_�ć^G��9re�K��I�u�*X��� (�
�v[��5c����"�~؃�����d�}*T�CD/8����7g��`��\���"�/ڒ�o��$��x�����*4Ũ����9Л��)�ރ �Z���v·�WR�B����}hN���r�II�"�����!��H9��4����=�k���7W�#P;�V��4y������G�U�d�厸'�zEL��V�b�?����/��{p� �jjf/%����X�(�O�~֢3�Ԍx�P�͢MD� O���"1�hGzD,��&ɺ	���td�Z H��A�ɡ	k�; ,d�U[[��E�_! O�|�d�҂Q���]�����b�ցBe��!00)�W�[�jf�i�^u�>�(�C���!*�L�^��H�yײ�%w�Xϊx�ug��z~K�ݚ\�����ib��R1�\��
H�f(#�Z�� ŏ��ԁ
$���ǌ�*P���7K��%�#�K�we`Q^	qv��E�����C�/��gf��b�/�T׼h�X���2P�ѹ�2䛟�C%~�:TD$�ԡ���G������5�ZI�����d�M��i&��b�L[L���4O�f�0�o�"�x}-"�&��DF�w[ca�յt�"*�d�Fjs�C#��7գF!5��;u�M���̛6JzO
`j��dv��z�������;��}C,Y2J�E��hP�B�9oh�c�@G���,��i_X������cm��İ�Ի�R4�����&�c��0=}aq�� �X�J�1�����|x�����
%�TgN2�����z4�X������Hl�t�p�';��ٝ6��+Djr��uW�Ж����U^���<׏K�^2&���Єy��x8��(nh�;[�@�=���pr�Q�Y{��v�q�K����ˎ5�V�a)�G����w��_,�M��Q[t�1"�u�m��8Vۿ4�$ f����}[�x�j5R7m�n��L�4++s�ݯ��N4fDph�|qa�����k�vf�}��ÿ%o���-W�s��2m얱�9���zY&�~Nu-c`P&7{��Z��
�xʯd]�M��g��G���о��	���_Ʃ�#��@f��C��z�UK���{�)��].�Y��C�=[Z0�/����e>��(���%+��	�2%�z�<>�Tz�𔺖�F�}��!<��<PD�s����lPc��6b]ӈ�ݭa/w�V�kn�������  ��`�����ub~&%�E��1�2�;ab7��������a\o�یI��zH�0u��x������l��]0��"�%�-���oTO�m3��4�����$�	�O�^�D��J�n�	���~{����`p���6ZЄ�w�D=%�@�bte��Z�ժty�.�����㨴P,�����}��-Y�d_��Z<,i*�����~Ĝ��� �ࠅ08���B�Z>fw�KYG=;[g��׭��mj%�1��׈<��X��>�����9n���>�6��d�
}2�O*�R�#\��YΗ��Ж��ݲ�`S�/<��%�:�o�.�j��R�������@��2�5�>o���FY��X!ۼ!�.8�B��J�Hw{�J_�B��dFp�H� CW����|@��W�ӔOr��}�p�h��A�V�P��j�����D����ܥ,�12SY�6��uW�xU�,��_|��1��~h+�ļo�y�
�]j���;�t+�e� =$��m_M��D��:�SV?jI�1GC4z5:ach���Q#�GE:�K����k?a=��;}��]���G\��\��n�d��Z�<��D�Hf�i��dε�Ӧ�y�;<�$�'`ǌ�e�V���G��ަ��k���1St'�ٳN$�0� �+����}�)Ӹ�A���?���=G�� �-��Ӻ� g��t�	���ĵv��{HOJ�k�Nf3>���S��J��Fiy��6�s?:�D��~�f.i��Z��P=mw�������H�I�n�/�z \�������q���9$:��*Ϟ��S3�>��0�l��Z`�S�'[0��E,u����P�#_����kqCl�r�;5=�O7?Xp��<%�"�H����?�.��V����x�Gs���$Q��5��^h��I �o��1���B58�n�bP�T]S�zy��8���y�5i눱�1F%��@B������*v�*�V��K�+vUm�Zi)auf8��'���H�B"��x꧗%����7�����2�K�M�,�`��� �j/�&��L39�m �R�5�Ѳl�~�O]�P���0��J�>؄���kk���_��Y����A(*]�e-(��ء���|Y�h��h?�M���*��Ew���	f�������O�&63M�sUj�`��s�g]��^F�\Z)���
��^��¹���X��0]����ͷ{
��6�0�^a�\��0:� Y�RA,���qW����+��>`؛n%�w�s
0�u�y���`E�X�"����
��_Xڧg�<����}�h��%$E�w)*So�����M��0@��a�_�ǃ_Ij�q����� ��[�v~L��ѕ0Wyk��{�� ���.��h�B�����ʢ,Eq�_��iDv0k�%�ϯ�S>�}��������==$���2%\�rGaZC�J>T�f�=y̝�����c��`��&t�&�����D��h�w��hvjZ�9�/y��/ԋiw3�{���D�l�;:F��U�ȬA(20�8k��������Z��TX�F�C"��f��ʧ9wz�{Y�J�-ȉhн#v����	���r�%�;T�P�!;��ݤ��
��_�C�I��q��YN}�E��N�Ձ���p�؟p��fT�6A�c��3�z�j}ޡ ����.6�����b��E(���v�/�VB�D���y�jɹ��Q8�j�=�G�m��h䨶e��?BfSP�"����xU�N�ʦh�^}zW*����1Ayh�Z��q����û}�`p �[d=��'�V���j������)�]]�G�I�F�g��o�D�!��~񗶈�lǭ�����O�k�^��q����lw#t����Mw���臱;ģU�{3�������؀�J38Q�e��ܭE���3�S����-�W	�S(��d��g?_�2�x�֟z���e&J�~|q��Nxyf7�L������Κ��։����{d$�#ɥX$��%�P�����
���M����:\�u�D�p\�@�*�>�܋��KoGu��o����8U�7�7�&KѤ@	�h_�Eaj�"��Crz��c=6���
�"uZ��۫>��j7�Y0ǻr!t�j�7R�a�nү{jOy�*�$L�.�Ye���:s�D��&��i���F�Ea��to][�^p$pl���zΛo1�i��N�H�`+�����̵��pa�**J�	h��ǘ"��Bg�MN3�ZKY�v�҇M�	���!3���F�Ux��o�q��o�_#X�3<��`��2�X&��\t��R����<?H?k>{$��W������t����[�HhN�1\�Y��Z�1�[�Y��x�@�����
����{庼[?��E�/o�̈́0��ƛ<�_(�e$9��&�d=�fܖ�=���7%ȹI(�{���R5����������? q/0L���-0��7�7?'�%
�3�i@ ����^$K[���c���st�=�
���.N��V�]qG�Z���>����~g�O�Hb}�_t]y�3�a�p�ʒ�����^��'�:3�mx�5�17L���_ķ���M��y��	����}��������Ej�t`uٗ�{�B���s_�S��$EK��|�^J6���w���E1�ݺ���wY��
��.�Y��1~�VA�y�[E�J<��Q�H`A��\�J_i3;����=�V?SP��W�v�DAc�����[���9��^%Yh��ۼ#{�`܏�T�#ˉw�p!���+!��.������|?������=[���G�Ce~R`UB�*�������<Fl b����VĬKH��c�%��PY�k���<?�y�Fމ{#��x�%	̍��R��1����{�]\Hm(�x[�b�wLW�aַ�:�l��*)�B�_o7��˳�����PWm�-3�y��8������f�����K���b��M��Mm�Y�V�KR�1P*P���R�+#2$xf�g%;)�@:ן�@'8 �|V��*�#,��D;5�_<��7�ӏ���)���A1]�5Ϣ[à4#eI�r�+�e�v��}3Le�t�QN��@�9��b��kW?��'�U>�6!���TTJ#����Rӱ�`������0ҩ�&R]F����V���麢|��=/Ǹ\�����(
}�@o|Y�F����R���:Ta�S�5���h��2�@��E������ L�)�G8�0�\���|�sc�ӫ�9��>Pw��{C�CGW�N}Ϻ�{�}�܁��?V����T}���
$��Euy�y���tx<������X���u�ͽ�c�^���6�d
?b+5�n�Pǳ��#97��-=�q�l,Vx��yd�{_�9��jM4��� �6
K~�Y&���_����  *������N��q�j�&�^?a5����Ļ���Һǯ��KX��Ik�v��S����b�����C��y��
�`��)Oa��E��&��)�J�%j�]FwS �8\/,�����`���\���A�A)$,�zmN�l�+�#���{b����Kx	1T1�"
�qP�|�)��!����.�<�������/Y�+�*�o�.�E?JOZ86��cR��S�%���+��}2�j���$�� �3 �����3����>����F���r@�*���-Pn蠅���ۭ5/��EPN��E�"�}��#�li�N>Q��1ȅۡ������>\�r4���>$º�uK�'����mH�_�� �M���30=��vE�XP,�="a"����K!*[x��M�����Az����E-}�&��y�ڦN��Cj�e.�>��ʩ����*�q�'B�%�j酹��[�Wo9�%��O�Q�0iq��ѩ��ގ�;��!����[���o���eMj�K����_&�?�N���|a���dgC�{ܯ�ɳ�Q9��\�i#Z��DwZ7��=~tY\�/7�NB݃6�4�{YN�����n~���.�`J�ހ�����Y�ҿ�]� J���BW�?����_�Q�Z�UF��E�ݻ� �B�ܑ��AP�ʹ[��GaR.F��pI�\��S�'��;1�� of�Of<5U��qyO;�c�~�/�[��)!�	�L�R��:kU���R&�A��2�-�������n��X.��0��U1�huY�n���F�WB���2@�HĿ�+&����f�fs�܅ؘ�g�rhƟ&�f��h�e<㛒������Z �a�
y�OR�*O���/A�|����'��܇�/�z'�li�g{���]�d�}!���-��mdH]	��瓱
�O�d�����&����_��(qy%k����WÚ���7��s�5^�PϏ%<�g�p�	���J�"�}�}Xk�b|zװ &i��*�%LZ��w�;I-J��?���1��R���ͫ5�`�:�~E�p5#����p�b�/Ɂs�b�+N��<ؔ�]��f��/�/�AX���J%? w7SЇ-F �����n�Гf+��]�✝vj�c��1ӓ�F��m�y8�I%T�����ks�Y�n%#��nb�*Hi0[�
��dB����mz�%�Ys=W��-=��u�.��=�G�DSkuT��
l	x�� r����+Q�xN/�~�d�0���Χ��J�̠K��_o��-�mf���H�Z@(���{�����N�F�Ug$�\�����:>v:ȋ[�jcg�Ca-V��|���t8�_���	����r�߿֠�61�ľ�roc��i�T\��f��U�]"s���S^H�Qp��*�&�ʋ.Oȫ��K�.�P��<�Wx���X�~<��pc6 _->�����W�lO����'F?�֒ק�l0�U��P��E�0�W��(�� [G;ӅR�I��j=t�s�O��
���D�ǘ;�ܲ��..Y�V�@f�~�Ҋ�)Ȱ��0���?�֦~Sx9��w�_����ѕ�2p�.�Cd%y`��G�R��^[PUy�pG�8slx
(t�H�����D[��.��(���M��l�݋�BY�Jk��s{�TdU�p�V�$��F�b�U3Ӝ{oE*s�F>�Ǐj
K"�	��#��L���:	����Y��vկ^"�o��J���V�l���CL�?DlD�zb��W)�<i_f�A����=)�Ao}F��v�%w�Y��fuM�A����Erv�37X��H
��z<򅘥��-������n[Iu��l�y��ϰ������"(��΍�ć�XX8�c�Cfr��IύlQwm ����wQ�Iɦ	���N�����k�z���M|�� ��k�r,���
�zb��:�u��@�b�r���Η�L+"�1���Y�"��kF�A1�n�:��ē�殼S@L���O�O���DNOԹ�	+����z���[�) ?����쳅�����+��X����I6��er��`3AJ�<\�M�(�%��Q����R<��t-��� h|ɟut��*��BzZ�����^;��%dl����2�):��r� p^t�wN�U��ӶAO�,��g��ZÍ��cG��.t&�����i_O�u��Z�.j���ONO�\�aUrBr!�rGid��q/g��~��/td]�`r*mE��do�d_b~�`��H�h�5�e䐂��|?}�5�Chb�3��;�qt���v_�K��"�o2jOM�d|42�I'�ɡDv���0��ǜ���E~\�t���.��>��,�lE�j�l�Er��5%Pz���-qI��u��.}�#&
�X�U�}>L�#���!�7&y��s1"���*|4�庼��Z�o��'C�����tJa�^�E���|���m��*�A��z�Mi����J'L��tk�X�\��Zyu�:խ�V�&9��>�|����xpŒ�QC�q�O}^l��E�f76g���:A��l#�N��˟(�R�f���; Yhn�8���O���B����O��ZH�p�j�6;ړ� I���c{��Ê`7kD��O�'���w�z�8����c5��R�e.��/��<��)ڛ<���~�ԧ��"o�CEE�w�q�lٱ?F��c�����^!�H��&���I��e��c#؏���!�ɍ������c�$�{�)`F���5�`�����e>��pC7�SY+�����)SB:����~2��4�����2���؋��3V��	;/6e�@,ZHÊ�V f�M��aF��d�KqhL�	Fڈ@y�:奲"�4���_�{9/m�oe�	$��F6�Ӫ��y���r�ep�A\�c�s��d���X��h��1�X/�����P��r����iE��H��έ�n������od��+���D���Cd�((o�˦>@F�t��H���ޮ��흪���@��R�E}�v�8C	s�^_H%&���cA����*C Tq�c%_`{_L�C�E ��Ns��п��?�q�7��"��{���R�T�m�¼(Mz6�fJ��R����ֈ����)�¯*^nZDe�e�/��7gf�)Y��񗲙^�p������a*�.Lܚ�Ѡ6ǊB�r�P���@��{�s�	���Y�cR,ޯQ)�%.�H���u�
�.�� ������c���x`��*�7'PH�~E���,�r����Ҳ�2R������b�7rc�ɦ���k����Z�w���#��d��-��ؓr�
�_�R�L��±�P�XS��T 
N�����tQ�ι0�w��I�	y4n�M!W�(���
0e�}Q�Djenl����)��;a�ɪ� |'p�^��O�?�w�[;��TT� 6�;@爰�G#ޥ�ޜ!�����'������&sw�.���WX7X^�@��qJ<ڇH���o��b+O�\ �2�:���ps6?B�KjR�n�,���0�����V����ׄ�����{�ܼp�F�D`T6��d;��4FE�-�:�/�J�(9�����b�����a�-AkK:ʄ�p[����9�@k�-ot.��f��A���S"v���#/؏,WC��+eX�wfq��SȘhY2��;OF[���G���&�?�p
��{��C���`[�VQM�"�Ѓ ��Ͷ����!ܧՕ��=1�i�Q���;�-@i�-�}zlM��!V5SD��{��fxYv딬����¦cDEzTj�A�%OJE7�B;�Z���c��r[�XՖ�A���9����C��=G�Zt���|��n���b�������'�t�ݡZPc˟��C�b��3\2�5@I� ���fn�H�������!��"��z��X�5���>����c.!�1��;ź�vyjf�&y�ɇ���RS�~���(��������Q�qE�e8	��d��c�\��R1��,F�O��[+�a{0=�0,E�L�����!���T��i���i�s/]J¿>�,��H.���6��#s�PeT���r��u7�QB��m�<��dJ��`����*��v��I�I��-��<-e��¶��t�6�(�0�}��Ys���mY�_1U�$��G` �; ��8|�Ig1�4����z �ÑZ��@�S�n|6Cn΄�aEE�maG��y�5P״��UX�1W�2&a�5�-�d(hK7z�����
�UZgf8Y����NM��W����[&�����cb�Z	/k�e^>�&�"9�����|(Et���X�e�	' �r"C��g��#S��|��{�L�%�����m[榆vX�QO�"kϥGpݸᵒB�e��D�{-�d���*#:��aO���mg|��F��
~���ꂇ:�s�8�^�GB��3�tNe}�i)�~^Bʀ�����v�z��-#Yi�0���UR��T�oW���
+�&5��u�;&]??���]���Ik!�ݵy��u�;���F�3`� �h82F4�u,)��=z�͖�oYx3n� S�+y�ǥ�*q)�����/��v����+��8���g�)�"�	�b�?t��ů�+.�J���C���v�1��Ǎ�rO]8�RP��;��"���&��eϥZD"+��N��6u��	���Ok�2;�����e4d�l��`VV,���	�U�C�K�\�N�P�Cc�I<b~|��-]� Ϋ�f��9B��E���݇K�u��0�Xh{G#�ִ�f�NԒ0o��� r�tI�	���ƜJk����T�9�}������(y?��7pZMt��	;���~�`�C�q� $�����N�=�D��cG�A����@�Z�N4�	$cʴ���zpϸ��T|��涾;�{�czn���3���ͧp�_���V��k_�+�>G�3�N�)� ?+"s`�Y��QwK������V�I���)뤇�|���} �W	����j�۱�^��àZ�㐊�f:MtV�h�e���O7�lX'�M�lC�����N3͙��<�I|�<�G�{&���� {\F��m���0�P'�����:m�#��B燰�>��aG �r���ZH��4�ê�*�8���AG���)HC?̂q0D�N����t���v�|7k�~�3ˮԟ��qa4+�ؗ:�g(�z��+B�(9RØ���U�e��~�q��
b�:�Q��(^Y|����+��f-g����>���r�����5�򸸽{���>�UҋzW�~��J��_wb���4Xτ�`��M���!^&����pl/���1��4�Aa SNw#�^�����Ӯ��Β���HFT�������Jr?��q�ʺU���(�ނ��ܳ���R����aQ�m�L���:���B��[��|��Ŧt19�|z��~Pg96xz8nB-�m���#Xi���.��|��O����̧���i$��h0�`������a�
Mxy �{?��,��Ch�J:hz���t�r�*�����!G��Q�5�̬=��pPL��v ��)y���`#W�U�U������x$���&����.9CphzV8k�b�9H�Y���^_��wU�G�d	č��	>��E~�uz�Jt����1��r��i�K�`�ؿ�?G�s�{
��<���.-@8Qfѻ����:��	�"�����a7����Ɨ��Jig!G��y�����k�Q1I�EkA�w?������P�AM�6å�v���iŮ���:��|q�������m��:{g�RC��;��`X���,n�V�&ƀ��-@�2�������Hyȅ�#-Q���dE�ˠ�MC��L0y�ߡ�+�J�Y�7O�7�R<������q������'by8�y���G����w���y��\��ʏ�c�;LS#/R��e�"� pZʔGr%m X������k̳�-�s��s�,]y��76)3��LuUziF!15�#n����X�N� ��
��ޫ�_U���Y����4������T�Sk&F��?2:v(�i�|��W�9�����Z�6�S���-1�H�����j�1��KW9�<cr紻�l4U�܇rc{����s�%%�˷�9��C�-�I�|�A��m�L6���d�{�}������{�i�f0��H�A$r�@�5�h9��YH�d������H�&��7��M.{o�������j��%NܗA�9o�T�j��JM��c�;A�ס >��b�dPûC�};FE���4Xܘ�պ_��[��)�\�>ym�\#���u(MbaY�Q��i��[ϒ"+sĻ�2�֤j�K�-� ���ȧ�����,�~z��>ʯ2_�K����o\Vb�mEę�"�B	�x�O~��+�Fz!�Rū��ɟ����LP�/�!�+vNgS�%�0��Le.�*0аj^;,Q�6*�r$�L�>V0��2���_�wJ�A��u� ���f�%�U��="^It�s�&�EF&�(M������'�C�O��t�kߟ�Wn	��U�m\9FuY�.w�tz=��~�GhF�\=s�:��yH_��U?�Y����ug"��õ���vCa�m&޻y@��l�Ӳ ��Ҝ/8�Hy�7��rV�����a�t�"-���C1eq�uU��p=��U�NR��|u�U��A�rl�,��x*Xf2�{24��]�C|�8��KȪ��L�.�%i����gљ����,��w8O�.:MU�������L�m�F���W�;y�ǇS!=lQCQJ䔝a`3M%��h&�-s)g!�$_� ��uJ�Z"A��8!�� L�)uݔl-�;��1;�lxu�-�Ls�|sR��	P6�>`��
}�>��J�E(�;��!�q��VV��M�]���ӥ������'�m���v�cQ�����BO�B�Q��HU���,߳4t��S���Z[evIP��������M/ՐB��{Q�a&�>6�HS8�XMsZd6NKIU�,
�S~?<�\�r������%=�%�AL�G��1P:������!�J���p��]ڀ�W����QBW���+�OD&���D!���}i,���b�tH�"*�p�l���y�ur��9����[�^?�At�d����t�q�A������Kv�<X�����jV����m�{˳��=����t�e�ż~�n����"W U���I�tM�U ��Y�*��P�QC��\�r�F��ex�Ks���a�a�G&��{�멈�6���g��)e�b��Ȕ;t
�:���f�m�Jn�E�M�B��o�8$���;[�J��tˬ�A�YXռ��C��Q��76�����f��M�V��Ķ�ր�ȗ�>�7��2���W}h:���9v"���mc�I�S��:/�N�j���>�.����Uq��������Q��Fbw��SJU�N�g��%�֑X'OO�j�BZټ<}r�)*�vB�X���7MJ������g�ϼ�lG��a���C�޹[F6�Β�%i��cwQ��W���<��Ƌ�=�Ky�So[�)��hDp���v�j��7��`����/>���r��ؐ�t�`�� �ބ.{����ƥ4?
w4q��l��L�t	t�@�C���`޸�>�6�Ц�q�����e�Jk~"	���Qr�����.�9k��eۏ¡�Z�7+돞����e_����`�	9�Y�̄��+V_@2{���,!}T��TxC�e݊��hd���Es�k<��/X$�jܺ|0�2�9��Ri~�����٤��k,z�NuiFN`N�'!;����Q.b����@�O=����]xP9�u�B���
(ֶ��	���Ed��@U���J	,��b�utJ6�j�`_�QBdD�]�����`lA`۾Z��Zr�M��_�%B̍b��x�p-M���W��'T�8��>�_�b�C�'_(��1��<�םPe@�1���@%:Y��ܟ�@��U��7E܊�.$n����k �2��qJ�OV�d~Խ}�*2U=޼�0�2���XV�����?L�/��lR��25r��d��7����k���+��,%qΝH� lۘ.�,>ͣ�dgz+�������D�����(i�<7Y��O��&�3LF��T�r.#�y�n��Tz�:��*A<�����D�a��K���{4��4)��;�oG1��0�	S���G"K�����������5U𴳁>�2�8�ׁҾ�.ϼ.�ä{0�Q���XXD���ݢJ�(�0O�"�w@�贈�!e���)=oˀ����N�٣���"=�+�N:��	���L���Z+��YF�-��1����nf���~�q�@Y	�E�x��'rJ��q�l�x�@�
Ĝ��ZH��p��d�W(p
��.cd��\1˓C��5�DJ�
�_���Z#�r��ϐ�rc�Z"��醝�5W|��,�y�V��LQ�'F�o?�-(�}4'3�4,(��mM������������*,~:#���p����f�;��>�}�[�J���`w!�J:j�)_���ZXtk��p�d����Bf��!���gVzà�6Z��fK��M^@e�W���lo,R��9��;�(&�je��D��k_$u�wUHo��2�����>��X�f��i�=���!��vI�Ȏ�UTM�O��*]f��T|Ӣg 'a2ſ�E[�G���Ϛ�2�c�I�)�i4��6Ԥ�ͨ��'j�>j ��uQ��xc>oW0�@6�j�pG=���uq�EYW6��T�f~�`��m~�0y��"ܥ�3*-{����&��ѩq���|t����d�=f�};���j�]Z����}���ө�b����m�hUlU��{z����U�j׌lP𶖄~.R�������e���Y\C��ޫU��X.!�V�I�f��@W��-��E�� ֊�5
^_��8��UQ��?[��H�� ��#�eZ�����+fgw\�L��E^�O�}F̌'�l����r��z%�^S��2�&��n�	l�Ҙ4��
�z���ܑ�po���m�h����*O>i�`���ʨ3��Q��Ϗ_�J[�rk�������3�??5�%P�n�����R����YFRUv
K�cE��.�@���9T��-{��n�
�,�42u\W���2�̥���G8?���kR,(����2��J���7��u��h�;0`�zD�s��H��N2������&n�*7��;�Q_2�>�JF� �6TA@��&8��rg^���M���d>QE��7��A��
GĻ�˹�s�ܬJ6�̥���o�{{p[��x�W��Q]������)��-��Ӫ{�8�ݑtc,,́;�m�����8�+g�� wB��a�Y�锋���� f+���!����D�à����������vZ���8IAH�%���S�N"�W��e?�-lN����v������W��럢�SFvx	%A��e��Q������T�;<U �����0�˿�B]��c�O0l[a����r��sɜ0ݯHʿ"h7Ʈ=��w	��3����:N�e0���-������iF�5���c�`���ʀ�H�xE��d�D�ol6���^Gl$�=rj�t��D^�:Ĳu '"�-3�����	r�Πy8c�A��pq̫gW0���I>)ì7M�(�؅�n����&���O\bU��S����������n�d�&Č�ni:'��(<�����ٵ�a�^����Xy^q�C�r�^��HA%�������}X����qQf�XD}�����s0,x)���n�[5?�w9��#;�~Vi�c�a�*��Ձ��i��x�H�'e궻�����5��h��H>��F����F��!��l�_��FzCZl���q�~�]hV�?� �:��\��e�®GuΑD����8�ɴX���p��Z������W4E✏ju��Es��:^a*�)S�3a7P�
��Sڞz���\r[Y����b���p��m�����)�c����+��H-L�и���^1'>�]dc��,�����}�u�|Ȓ���ZH4g�1��X�2��t��u�+�p�^��	�����?p��I�Vq^�����:?wJ�;DsO�Z6(v�E�.�K�&;��`6���þ�E�'	�{[���xiM����l�c�B��n�}(��4=��
L,�����Dy����(lSe|��~�����V��fp:��"���h�#��mnv2�q
Z:�,m��%1�&�+t*��#k����{�!����f��]M��
�z����p2���B��KV���s=i�2��xҒ:�qA��hc���|���O̠/m1%$z���$�};M�`@��%�Q_�wÚA>�5���Ԇ�@�)	t�j��(t�PL��q1=�����:DX_�8�7b�C��K�j�Z��EAf6|�%f�Tr����l` �H�s�½�Gx��5^����yz��$�\ѧ�g',���������F�,1����2�Q��lǤ�b|�7�N��'1-����q�X7y���so=zr�N CB��L����S`�3܁��ց3V��T��2�!��:�c��^z�AGX�1��B�4��V�+ox�Z_S@gӭq�V��$I _�<)V��I�%�H�%�����X]���:s����X���.�Dy�N՜�5��}�%�5 ?S �����	�):����ANŉ�����
�������6�Ն��h���תk�g�m���-9p��2����汉����X ��Hi�7�`���涿�F$�Z�����K���Y3�u��1�.����'�#:���)(*G�j�fd@h��Fχ���g�~ă	�m��ɆPLs^��8J�R���kc�Msn㐉���k�24YZ�hy��H��kk����S��,��ހ�~���A��r��m�(��V�Pjߔ,�����ONH��b��T�F�Oҵ��� U}	�T�h� |��;�����X�^[q[��@�Oj�����O�(������[�����������'^S�.�Xh��$Ԩ����7}�>����D*��Y��&�%ă���bv��>tl٪�]qV#���� ���.p�P�`����:���$Sm��y��&��6��`vӰ�D���W"JJ-3PtS5��b��n����r�\9Mk�oǐ��r�L�)񚡳�ī�%Ǭe����i˺5��m�"P7�Ek{Y��E���#ʻ"S���D&����Y���}y��4�ٍ�+�P��U��R��)����輇�VG���n��� ����������� ��x7h򇚚�zg��l0��tS�qs�K�z����	�����yCv�m�E�V��El,�J�0z �C���ٞu�����f�lX@F��	���\`�;��͎1K�J�m�Oj��U��ێ�m(��~��H�4���v�Ӿe*�����*���K�#�	4[�?��Q�����{3��Wޡ�S�2ͯ����p(���h��d�D_�En�_�bwΆ��W8��ݲ�p�����x"�Lz	� x����9�3��2��Ul J��mx�J�cVް���4|�S��L�#ش�ڬ(����ݚ������s��bP�FT�հ%e����:0�Od"�-��;͛�u�O5'���&��J�L53M�Ҫ��*�MR��mLc�ј��|�SZ���� Pל�<u�#y�����o/��
x�Tw����#��ELBOb�x�����4���DT���6m_�l�ǔ�i]�(X� f���P	Gj�w�̺b���i�.ƥ@t�Qp��c������8�A����L����SdeQ\�&0[J��Յ�Qp��-w" m�WY�^G^�~E��- x���x% ��85�3!�M�K�B�B�9��+�SB]����K��k�Gi=�K�ϕ��-�ϛ5��|������s �j�(�~��Ln)i��E&�����^���_8�z�P\��Jʀ���މ�Ɗ�����m��r7 ��?%#��^Ng�.Ng�|�B����9�����AbX4��\d�����\�V�6}�(���ˈ��<�y�n�r��ت��_��y� I*~.�^���B�:+X�x��[��G�����#WO��:�$ϭϒ���厝0�����qay�(����[Z)��n���G�\�����y�+�W�4H�=��	���VCk���TVM��b"l:%�vm'u�e ���
��]�ĖL�����Hĭ֓��yQ=���r<�b��&$|�|��e.(ͬ��7�m~�������7���9��x�fC��$`�Ja�4���Lf�Y�w'\�ʇ���A��K���>��O�@����+	V�z"������o��#��1^g�"Io���}bϞ`7\�<| D`x礀��9T�q�4�e�$�t�����q9�ٍS�^���B!�B�	�Ѹdބ�&7�sQj��%!�p�qX�f<a�(�8�͂#¡�|�E�*���w���u�v��z/u_(�z2�:d�#�u���D�[I���Q�/]p���"S�9������{'i�Z�50A��Eh��Jn�Ed��~fi��������S��y�z�d`�<�����D�:*��6��r�"�1l�]z���c��nF+���H�Ԓ�=�h4 �9�'�W�7��:[��]��yh�h�7|G�~3����kA�P��-�_�"�nrםv����p�'���L����zez�_9���u��B7�u�;44�xL>��^���EH�ă���	���'��X��R��0;����J&�/e>�i@�d��I1_�x��d*�Jﹽ���Nf��(�r5C�$����n��6�$�cY�	���
��B�g80�����U��P��a��V��:����k�	f��I�~*6�2�P��|�9+��=�{(��6!{��ɺ��H�'��}9��.^X�(\�İ'k��l�RWq~���(��~�������>ȡ�q���,�s9����x���B�1�C��w�¸I����=C����(=&=���:E`[Y��b�J�� 	r��W� �H��
�T�+�2'�ܫU�T�����^��x��q����r7����2����x'@1r{���~#�3lD��+��ڵŻa����V2�a�WC��0��%H��Tmҋ�V��*�ch���U�����Ǝ�W�%4�֞>`�<]Zơq��Dc���Y+r�_�&!���ۓJ����n!��ԎOR��jPO�F�e�Ƀ����r�8B.ޏɀ"�e�ݠ����~�}���&�~�|�(vG���o(����=S�,,�n�!�"WU�Yo�h��R�~[�uQ��p�����؁��z�3�'�<S��n��PL�Д���R��,曦O�;�2tG�LY����*���p��i5G�O^Gf#gk�^y6�<h�^�Ìա�
��K��4$K�֓��Lj��$;=ZO���n���o7�>l/��;��Sĺ�����|N]��-p�m?��(l��K��w�X~Ԥaπ,�S��HE���:k�cPa�E�3��0󿸡��f��_���8%�_�~�8S?�s�޲�΄<}��k%�w*��l�I���aS9��t5����cҮs���c`.�uw���+��w�� e@7�d,�>�]g��2
��,�[3��/���AYٴ��g�j_����"�Ya���$�����3r�>sz⽐�0��W��D���-T�D�z�4�G�R���X������<πh�}�G;��i]����C��V� �[�W��S��[sx$�=ۮf#S�Z�K~��wED�D�x�{ܮ�bl�}��F�s.�e��bKN��Ȇ�<�&�\�&�bMO��?�g�� .ߥ�8�B���Qt��b�����]���؃P;pKs������!G$�s��k��l���^c*&h!��-�vPk��gN��b�1v��,5��\��U�H����ܔ~kh�X5q���9M A��5���׻��ݬ�̤�'�u*��S�d2�J)C�rP�?.�LΆ�$�͛�<��̼�	a��f'eB�H��h\�_�-�.Wa�E�aW{����=t��8ۚ��LcC�|�!�� �(��ᬍ�#$��~�=���>sQ\Ԁ��Ot(�[:`E�{֍�6��C���� a�k�zP��t;�mq��d��X�k��}	6f#�tf9~��|�Y�,<r���V��;�����j�O��ܝ�:ĲZa�k��E�^7Ry�T�6�V����<jWS�k���"��^<��w�n��&��2�z��.��l�S�q?~�-Xf���i��6,׈UZ
��J̼�Ծ_����e;�6�:y2���� ��N���.����j�+P����Y�5V�0/jG����� ����\+�7�9$�C\�1۷�ݺH����3=G�iMc� ��4�Bg!r�%�E�� ���z*��*��V�*+���Z��6��E�k�u V03����:��H猂X�3v�D�{3V�D��g̒Vi��D���CG����碩FԴ��؏�R�5�)u�luW����ђ4u�U�w�����ڜ�=��#���?d)�����;O�XCG2��v�$)��;k��3SL<1���QR�'�>J%bx,��V�PI�%�Ŀf��>��u�/_U�̈D�P���7�����ń�T��p7g��Nn*b�^BG���N3�-6�����_>j�P.@�����F����Fҝr�ӊ+r���hJ�?:ƚVZ+?YizZ�%f��Dп�R:i>�R]��y�P�G4tESJ*�8+��7�.	G�t�$���t��݈����V���q��{R�Tqn�3�9�h�^^�#���C5:厘�V|��?�_���649}���;�ﭟT�B��&��t�ͼf�z�Z�Y��O���}�j*�ڇ�4l���u��V� P�(;q?�{��zY	��r���m�Sn��'��G	�=�N�;������,N�	&F�: �j��@'.\Ԩ�h�_��ǕaGUb*�4����A(��Q��+���W~d_���]Bs�N��3Ah��|��K�Q��K��#��?j�0Al�@�P����;��	FO(�q��������y�
�!ν!k�r�?wPU<���3��`�=����vi��;=��p���w�I�3��J�i�7��W��>�1H���V�J��Y�a*x�x�>�9ɳ�D�-�Wy��	��YM����M�	��2Sq�i�G������P8�mZ��LB �G��mw�9�z�u�]Ѡ�֕����5G΅��?���M94ٲ���`�wn��.x�ヾ�!X�8�7poÑ���Pk���\8���(���bMT�6tTtpҲ��|�	�`����e!��?:v�����+�٭w�5@�;%Q��f>B��ֈ��#n�ut��޵�-(s��VN�<o��Q-?����E�M�����&2�lG�!I��5���e�፷G�;���TӉ�
���|fA�_K�^l�2�a���NY;k&��m���F��,��@�-����詪io���v\f?�>q���F�l���@�]H$�w��kzaS��z�������T{��K3� 2�d���cġ⍌CS����d�F��g�m@e��ܰ��ނU��-j��q��a2����4u>���i��!�y+�/*ŗA�؄O{���do�ip�;ZH�7�"����VB�D+���t`�7
��=v�q��G���cjcz����~�ᖽ
���1�$�a��# NJ~� �ق����	�(�/e�J{�O(�_�x3P���Cr��\yl�Jx��u��h�~�ׁ�G�����Ϸ��ׯ.�q�xx�JBF@���C�q� �Ux�~M�8��Xb�F�)`��6a�cݫ��5�L,�[�����d L�Ɋ_9����h�����+8@fu����y�n�n6�88�w�R���N���z�����3V�L��<_P%�Z��@���-�x
�n�ԅm�0�T=�$9ȋ��4	I-I.�t	~�[cg�ǡ��9���C/sB������L��}�5d3��i�T/p�-��M]�$�69��5��.� L�f����T` ^^�ŸЄ�S��z���y\).mq�~����a�g-@���/l�.T�Dv&S�6�D�,�z�U0�X}����(Jt6���V�,��]?����d����]iw�)��+Q�������5d����K�1!��tݶ���@)̦�˲M^� ޥ9�{n��0I�v>m��Z�����������Zj�tM�qU����b5�sp/G��$�s�l|��1䙿/���[����J�57e�j=s��:���2!�kO%�i�x"��Мj�V����\Ѱ`佺�GU�I���)ԙ*!���{�7��Ԝ~.���G�|J�D���,$�|ʂ���?�B�	��4�������g|%�Ѹaҽ��\�QC��詣�4��>�rK��y�g�(�����/+Ă�����S��G�eza%��r���x�|��&��)�������V�Dn;4���-OD��&>���s����h:"BV@����������m�,@uRF9��l����'�����rv*�	|;z*����P��q��҅����mﶀ�Viz0�sV�k����EzE�
��c�9�����@i<�VV��Ŕob��XMX.]��p$ n�q3V8�k���:�N�#sA����4�����߰0���f�|�.>�AY?쎣���Z�L�/�X�����t���S{YN�)��ެ�I��k�K��ٟLvru����T�|�V���� �6����&}[�6܋2[�!��Zgl��-��zF��$�ɥ����V����20��
;�O�:X��h�%�*���V�9�0:��1�����E	[{�I��%ޅ��5�ݕ{��*k-1��3�W�����
� ^p������Ӛ5yJ9�8-5�x�k�d�*+5Wb5f�N��~7 )�w�V`�h3�PYJp��D��H��@H�>�^� =U�D��q�y/�U����;4�W2�i)�469���5���% '��C}�.Fv��JG5/!��/n�N���Y���.\�ȁ�g�|z8���ώj��6L�wϕ��E��x�Y�Q+��'���H��:� �H�v�6��7פ5\��3�L)�q�w��bj3oL귊�����gj6�Z��
���gO$�9sp?R���W��1O��%c�q4Px���bjڣˡ�r�Ι��"�b��ߖR�a��]�K�b�L�qF���aJCMN11����1D+����jۡ��)N��Ip�<	W�%��L�i�[�Pzr������;B������G+�Y��Yq�mǞˬ=g��p+2�a$L3�e*�Ĉ�p1 T�QXz�r��H�!O���p��ʑ¸���m�^W��"uk}�iv�
b�w��/�����W��v�E0���W�DvS�����W#�c���x=���ȅ-`���/\�!�@g�{ծ���(�D��X����C�è`�G��Q?F�āw�Tyvz��D�e���h4�%��A���UE
y��aF^xf�3!˪隆�:��@�V� ��U�r��N�l�-Nb���q��k4�����k�p�����h����Ғ�-���M+1��T�d/~ā���-�fR3T��A(?ӱժ�Ԋ	�`��5�Fm�(�,DSv�G�E�\-�r��Hy~����n�XHOVY�μ}H�,u���ЁdUK�\|�.C�,䮒�e��7PD����_;���W��G��Q��$�q����s��rD3�#�����+?�܌��ſ덊(����fq��"�pʝ�+J|(���{��@37�Ř��/n�$;i��_E.��1X�g|iaU=����6pz����F��`^v�x�V`�[(��W�O���*'�HN8��)�Tx+J$���	>�|�D�Ås�p�#�@���^a�S&kf��[�oy���kxk���2;_��q�z�_9� 7�7�n<���W�\�0�C�*ڔY�vJC2aD5��w��fY���uk{���\�5"\�GD<���'g�+�a�� z}b� ���J�gtn{ӗ��pG|�ٻ�D�:r�BA�~H�c�/���4����
��@/�d�p��--���m�Kj�m�
Q��޵�
a���+�Uk�ϞDx�����}��}g�n��
�&j�o��ܩ��Np���1(�rZXv�c~���ƋGL^�ށ�l5s�X�j���EkCr��͝�Ʉ��Mj�P��
,�n�/��h��9��F{D�$*W1Ŕ�e��w"�t�4��;�k���l�V��l3L�&C������� <������O��>����Gm���L_��!`��{����W5࿋?��}o�pACDO���th"z�S�SO��[��$O��aR �_�%g�	fg�[;�'�W����7}�I��	��w�}XfBhie8����E�x�чe=�K�Ju�Cv�1ϧ�	�Us1k0 }h\������������+}#�v��\�&Vrp{����t�r�:���ZU_M�����V�"S��X,_�ۡ��VF.�F�5��h�t���Ñ%!����9CB��VH�o���``E�}����Q���1ԙ(n����0&丁� �Q)Q��1��pt�,�kG���:��O�B��n�=Xd|�������akY�+�<�����UӴ� w�UO`�����+瘬S����u�H��Le�ê�G��^�2���Sɇ���J��&/�;�{6i�� I�ܞ��%��_9g$z��}�������/�ka�3iT'������>����B���Ns��ȿ5�#���:�ūt�N{��k>ƾZY�g�m���h����$���{FO@$����nA����Bh F��4��[�@.����I��x�������Ě?c<�j������E���cֵ����k����`��Wt^`�͑_o���iT7±�i�&����Wi�Š"H	��-���=� ��i���iD.�'����*=7���W�V⟎-��IZ�������5<�˝�c�:�n)	�K�i�j��y�Ez�5�O�fV���W����� 7?�^�m)F#/�w'�i"�f��A=�j,���v����MQN���^��Vi��pg��y�#��[��>�؄��~�
��C:��|B�!RA�}l��|a\_����Y:UPW�}a���:�>�Y��U^�F .2�Tx���įÜ�J6�F�o'b����̎��p+N�S��s�a�D�"$�%췁��xv��sgTEz{��_U�K��;㔢��d���Z�X7H���-e�`����۵��X��ݍP��niU�x#�xy0��_��yW�wn9a�B�܄\,�u�LFYxN���gn��z��)��&FAZ�'�W�u�������Y�$[h7�<�[�P���E��ոuȯ nz�Nz&KJ��.ĎW����O��V+\�3>y2���k��ϪTb��Q���굍��zg�r�Ʌ9��ɯ׀X��b���ѡ�7s�7>�L��H���3�h�k���v� RI�)�Mw�/��T�{W�R�dc�?�lp���za�]��K��	Ǘ~2}�ك�R�8�\�b(.�X��\I��� )K�p����K#:~�Ń̝j�D�|��/�>�Y�B�CuTZukmMx3h��Nm�S�TG�^n�#��7���-aEj  �W�M�1�R�f�:�n[�Hl��o0�=����,�/�vr�$����pd�|�1�o���Cږ��m�?��3�EH���C��#�����U��ihO׉%#�5pY���qeLg�����J�_|G��%�k�NI��R;�T\�� ��LW���mu�#��6 ��h���� ���-������\�li�����1���������<��7/��`��<����l���ש1�����������Z��¡�P(�znx��H����!J]g���żՋh��`W���?+�B=��}�4K�XV��+p��'dl����\k��L8��F~�A.�ϝQ$���29�t筽��Z��+TK��GP�G�W�T����c�=����!	���t�sd
� L}jC���@8$���W+�{�:��,V���EnHI�L:�~��T�����#Z�l�CT/��L`@�T����ǂ�U9~��Ǔ*ab!���O�)����O���u3�dt�"`��p[n?gE�O3d��(�{[0~�?n�%�*��LT���:���G�)Rsx��_p ��$��&���o�[��>z�uMl]i��t{ ���(]Wǂ;/����R��O��o=��}+39�n��p�:���T�� ^I**�ט�Cs�����`�]2q�s������q����L�(��o,֨|Tэ$�W31�:��h)TI\�;�zҨ3lv|B������5U�3�a���:��0�ʗ�r8|7�����ͳ���@uQ���<V��v�jD@@rXʵ�5��L���i�B:E�[~���L!e��ļK��ˮ�o�)-k8s�b!l8�.�(L@�;�p��iE�IEnY��Θ�h9<��C�Y����b���⻿���,�tWq��zHb��3����H�Em�}=�ݡdt�����)���l��հ��9�}�JJ�A��ì[��3],��ğe�t�ǻ�#�E��7Wm�T��Z?���t4P���yl��I35Q#���,��*W�A�6a�s���"mܙ�W$YY��1�hx%��F§�o�����*�a��w�XV'�'��E4^�h�k�?.Z���OgI�2�͂�|J>8�0���b3����#��\�L�`ӱ���H��
�%�O���vP\����6{�X¯n?=�n������D�S�����g�|�=�=f�'y��m�h�N��R���<Dm��Qr������`����,#� {����,/���7}<q#�Y`d�%��L c4J��	a+Fo�D��X�ё��r/6>��KFߜ��n�^�BOFYz�:\b�*��w�>��2��qԘK���:�sA�j�Vi�M�	+y�}2fz_��jC�l��d�gS+QV��K�S|�h�Vϡ;�ǭ�P�_~UÇ�4u�&ue����{/ʳ�Ll,�-Ba�8�Hw����[Y�%0�xS\��L/#9�3q��p5.��A&��H'��,^\_��˜��_Yj����f�Y����Z�S�y2�ZB�f=啈oTL��G�
ؘq����TT�c�ly}�H.Pt�	V�/ʴ��w82��F�����]�}�,���{ ��]9$�m�V��A#{!b�v��?�8��~y�>���'�{���Y[a���ɔ�D�-��?5�U��F��R����2d�J���\Q��M(A�\���C��{��FZ\g�<��&rj���R�B�.�^|QǕ�i�u?Se�K�Y���ss?7��6�Q���݀�M�Vz�3t���B���Pi�K��D�����w�`��MX̽9�v5ݹV�\l?'Ƈ��r��Qu�q,�$�H�s�\�YxK�O���8�fwE�>^B5�G_��U�ab}{4�f}�ɡz��}�.g��Q�*9Uv��Ź1�8?��<�)��A�u*��q��*ڑ:R!s�5祂�J�!>���C��}���%�����%��=C0v`��-�K�-��B�p&��+��î�;��B���Fa�1�L"IN��:��AЇ�9����IWW:)@��q3j�X Y�O-$�9o).k�z U���[B��B��>�Y���R-<��O�I I �1 �x�C,�<����_pڲ�����������md��n� &c�e� ���<4�����!�5M�q*	k�C)���E���҆��m(�Nm/ -�^KR?��Bf^��~,�W�}`����KڡJmN��Q�m��g6T43=�d�c�y:��i�������ys���kV��W�c�~-`�8�4:���F�u��G d���Im��D�v�i�ġC.��~^0���������_� u]8���..����r�*�)�����;`�ь��4z�jlB/�ȫ��[����jw����˯|L��u�6�_]T|�X͒�%?� Y����Յ��KŖ���O�MIM�O��e^nFݾ������+= �@t�jJ�V�1��=8j�c!�3.2��ec��̼ы��ӈ]������t��NVR�,*�u(�۪��7*/�21o%��d�M�E4���o�%��0���*K���FY0fS��c|�6�f��� I�3a;�A�Ȑ���%��!��&ޤ\��$��S|�/�3u_�a$簇b�0)�f3W"�ߍ����2���,2b��br%<���W���p]̲�U�7��ve��T_	,s���>�{���`����!\#?尤Y3���|CHY0�1�y�و)Q�m�Z��(�Q�#��&"������R	�
to~~�"�o�\���Ң�� ����h-L��~�`P��� ���i���R���P��;�ئ�f5��)��)���W6��񷀥�V�qH[�݄.�z�B�Lxq��b{Pj������u�����Z�����8��+x�q�l��mD�> ^"bs�����o�hzV��} W[�dKq��1��*��6D��7v�t��eD�����J���b�j�H(I,-[�R�A:$�u�B?h�/lk��]6{ȍf�����.0��t)�i��>���=lԁm�ф�^����=����`��}N��O�L^n;S=�g����7;���<
�D�Bᭀy>�C��������J��Am�[&#��G����>|��	�4�f�AB��Sɍ���dG�-�ۼ+�Z�J�>��x�W�J���#�<�V��_+�k�V��e���l���K�>+��Z����|"J��c��x/3(��l��R���6-��D0�@��E�!��)�"�aEKnq��r��%�Km�ϧ��e��rmC�#%����n��ӹ�'���R'b��-��w$ߏ�� ������*Ң!9,�ȣ1��F����8ӫ�'���¡����Â#�*�ݤ���>9]�h��^P뵘�4���c�>�|���Z�Ͳ���p���#i�h��R���{�[�3��e-~�ٟ�c���u�}@p僁��k�|�Q���y��ga�~���$Br*$0���b	�����klN��"�a������Wu�!
e�L�1`b�$���T.4[.��7>�]�e���5`��W�`���6�[�H-�0��f��I7}�L��WZ�S�	N�*I:��ݞu����_T��-|�_S�z��Lѻ��|NQ��$J �%?n��'��������B�2MҜ ������}PN�@�H�p3����_��z�k�kj�6R���g�է�K��oUS���3HUz	�+$4���=�4��� �XL�lESM�9ݜ9�As��@���[+k�؏"�Y@�d��כ���м�)���2��|� ����0���,���-t�;����+=[Kъ���U�h�q����F�
%��W�f$�;k{m�����ӯn]\ɺu���̤cf#���"��?~3�
�[���T��aߠV��L��E�.�iK�N��'>^e�q�ߤ$����@;�V|�	1l�]�Z���V*���gQ�b� ��Ja��-��D�N� �/Xa@���aMG>��/�j�0��0-r��9JCK&}�@~>���$���.��0�թ'&�OUz��\��V�XKH0T?AX��#��3��L�c����̬�'t�r��`'h۪K�~7
IB 6�����j�yr��3�\�q�����*4�w���o��5P�W0�[���<:�_�� O/�҄�5/�ޑj� E����Y/,�J
,����,���I���^�
w�I�
�������u�H�ea?�I�u��PF��t�cK�:�o^���7H�����bO��r�\eqf�(�؏r6�d1�P�Ǡ��Q亃�H뫪C� ����"�I�4x
Ĩ�m'?��U��T{vx3��o��N���&V�I����μA8�'~���@���"d�>�,Dr��(h�I�Nؐ-�i�i��_�*��ua��J1q�'aͲHɦ�8.L-�C�Þ�9�P�Â��ޱß�*�^59�����U����p.0�Ck��j5 ��:��7A����V�;)��Lv#�l2{�4��}��"�Wʇ�{|����Y�*�南3?����j1+�-�=O,T��"T7�=�)��,��(�H�U��Wtͨ(Čr�:�y� ��5?>H �x�B�h� r"�7���W�1�e����>5]�09@�*T4����w'AU�)����u/�9��Bb�?����O�18�����5~'Ɛ�9���&�GS�����A^���P�K*�}�s`�_m&�-^!̰�P��t���K[D�2"��a�3�����&oB�KH}��S�2���޹�p�D?����NO�^=~R�?J}��c�q��c�˞?�����t	$�`�V�%w�G������٘e��؍Iԥ�U7K��ra�@���a�86)�"�*2C U`C�1.�@�HLMmDGmL�R�P���:B'��B��o͓WBj�'�`�՞���O���O"���ۛC���D=Ͳ�y�.��ر����)��gm�v`6������GBϖ�˝��6�-�Գ��ʮw>��6�0)�\FG������v�y�c@��*'e@�ᐏ�`�3��}1�;�;�JS& Brs�[� xf�!�2�t�����l��^�N���?K�z"|��dy�;ܚ��`�ܤR �h��km�<�RP9���acFhy�R2^�?�P�
{<�
�g7��<��gK�p;��_�e�l�/��m1���1�	+ ���Y̅�����m{э�9�uo��*�	!wpwA�}d��+QU�^a
�b�Ov��o�5$̜V����:[[�|�|mYͽ��,ÕA(���2�b ]�~'%�������/5|^�?�0_5�A��,Rv�0t�T}�E��[��E��Ԙ�=#��*N~%=/WU�>`9 ���9x�w{��B�v}\݂{~M�#����^�"�eY��^�//Ti������� ��~rΡ9c��.�d@a@��5��h��DMETن2r��:RP���YgNQ7T�e�� ��֡ƺ�d�?����<+F���(L�i�[x̥x`��P��gG�T=E�G �N���l=��;�z�X�	�vȧ�޵ Z�Nw��{�[CĈ�ۨ7�|ġ����+�R�.��a���ҳ	�E���#W�&�12Qe':Ts����'cǛ��И��c��[9�L�?�si��<K�Z$��v�G#༹��r^Y�\ɝݱ��~��b2�P|t��IM���L�ډ��PJ
�㑇�~�P�>��wFaqYl�!*�q����`�ҡ�`RN�'^c�=)��/	��txſ+�0G!����d�����?.���h���}%���e��uawI��"5��n $�8	+Ȅ��_*���R�wkS��#�:����۹��y�߸1_�U��FZ�]��)o��ٻT�!	��GI�+�����Q�
G��n�Wd��km��[��H�G��nc;��l��| "�|�uԬ�S謗���^�5���Q��k�S�&�lh�o~����K��*�S�+'���A�"��H���
������f@��{�ǀ�5b��ȓ�����~W��R���[lH*M��e��Q7h�V6�{�(���Kr�ԡL"���%\b �I| �4��Z��� �k	�*�>-���[E��6���ۇ�I`iA����{�d�1��@�>Z�����J��*�jĜ`����pͭ֋�7�T=���޽߰�1��V�FE�8*fm+��$� �$�M�z����|,	��A�.}�+]T�l�(j��^�^4g�X��*�����|m����4,�a�Z��@ִL9��q�s��}�A�/����Bl��r��J>�_6�K
�@�Tu�?�	�PR`��q�*ߏ7��'x�mLIb�=̻�So3����"��>�S���_��6�N��'=��d�����2�03	�]�oQ_����z�Z����̢<�QP����?ӝ�z��	�}�# ,z��\-��*W��.?D
���8~�=!���ZљR��g4ڴ���^j'+�&�����?��y���_ ��$.�_�V�0��֬�e�údb�Aa�uNC���uۊ��Zr���v{7�L�z�H��S��(,,&9���AM�Y�̦���|��8V� ���.�ԉ�5�o�~��[`�x��$�+�%%T+�����/�.{-L)m����$Ǯ��b"�e	X��5gKS���|#��r���j4�W�&�k�p���D�u]Wa��լ���>#��Xkٷ{���$+��-��&& C�Ѿ�Ͷ��Դѣ0}U�f�R�2�py�ga�
�c�"C��F��G����,��Gh�������}��;Uũ+W�����B|6��A��{���&�DxN�q��1�Y��6 ��H.o'b������vo^��z(��Ks�Y.��Y2N
�Aj����Nlܴ��h��P�F�Tia>�Ґo®޽����Ԯ���Q��|�z͚;_�`��E��s|��to*���Í�b�\}�ك�궝�j����I���s8�(ǣ�qζ�@4*~䕵R��cE��F�]$����mS�rC"��y*^�yax��g����n�F�`4V�	��Q��ж
�О��ϝ����R��Hcg~�}�?kqpo'��!�$� Aއ!�u�VY|� G��ЙsE� ���|�Л@W���*����@�&s�R��x=��<a��~��A�����:�P#�!(��g���Ԯ�)�W�
����\���Z0�	����h,N��v�9��R5��u-{�+o�bDzv��p���DlzE_Ys�������e�>?2��iuL)츫�%���O�?M/d��W���^��3#�<w߿��͟4{z�`��҉�:�vz^G�կ���vh����W��%#
�e$77�sF| Gq>ZY~X:��)�#В�����m~��!�l��G�k��|C�H�cnIv��(�U�&����i�;&�Ûm��� f�C����F�a[]?��!ZC�P0�]M��.T-K���b���U�F\{H���״U��jǿm��V��	f���._{H�ف)p��P��Y���0��������	�8���ܿ��QA����w��kI�N%֊
�P�iW�G6yv�V������E�D�(x�'6�����x��E��ѡXu�56Ob�Վ��H��1�|#l*LK�Z~ͬ�����zy?��E~���(��p� E�m�;Q�u��H�ϊ�EΉ;�}���:��X=��c�۲1+Dk�T������ƴ�'To�0���dLa�F��:T}:;N_��K^WNF��K���֯��2擖Ϋ��������kC�� �5؉�4|��O-m�/*��E�L���F��G�s�ߊ'����J)U���D�l\kD���T�A!ӦZ�e�gN�i1�s�����:�M y�u�cԚ�t�1?2[-�ɹ�VVԁ"�KL;��y�4)����m��F�o+E��ĂJ��uƉtZ�qc���@<����p�����EFs��	�7����JS�ͽ��L��k0�8r�Y�+nd�
PѾ�*e��8�(/�r�3����ѭ��n����n̖S�
�(�
�Z�T�:�%EO$�(� z_�.���(w ��[w���P.EV���7+5����F��|��X/G�0݄]����K�����W7��<?k�O+�Ljs���������c�&�G+An��tx��L�)0`H��6BճBk����E��[�.����i�"H�#>��1i2O{�fP^��|l�S����o7��}-ꙣ/4;�@>�q�3ȏ� ��fcD@����mr*�,#b�*<��u0!���A7�P��4m�bȄ�7���,b4/���ׁ]����P�X�ٶ�(|{ӽ@�����B�14�m��8�_�����e<|��(�3�5z�˿y �)Ȇ�����Z�Ć�	����G��8Ca�r�(o���~hV��1)v3��tXrW��\�Z{���,�7�]p{���H����w��}P�	G�>�!�g����iw����ͨ��JF �V�0���i1d���{���R��qv�@���dt�1L�h??L�l��#�?��k���E�.���b)��H��!��nv �'zJ&݊U��5���b@��Ȭ�G;��.6��V��$S8�x�F�D�꫄�d��+-�5�X�#��������bt�}<!���h��'e����#���(��$<��բ�Wx� ��:Z-�I��ot!0��;�w�A��j�J�s#��~���<��,s=��]�^ϡ��N���r���>�w�ج��}D|Q�L&**�|�ܗ�@��@��3�?\�,����Nh��]`��b��T�w�N��&�7���r�eq���tK������,1��j�[�H���:�m�3`y���k���?�d���W���C�}�?AQ��T���1�%�~
��t=�O��ȶ��m�[��7�u੎{������ˁp�8h�	_:�&��w@:��\@T�G`�e�G�X��6]��kdM�tH�.���+�Db�P�18���rtVVѧ �<�� ��9�MX�D����c��I�C@G����o;Hёy����M�>�+Cl2���Fx�i�>�#�akK�>;��vnד'�졑+�UzY"��nsXn�����๻$���G�e�BUd��Uە�fI�{ ��gŕ6�k[<tx,�_�뺂�q���oGw<�qbF������]��tly��©��A�,�7&u�o/
p�H�U�?�5�}:�����b8u��^ScyAj?Y˴]�E#o����冤�F���	0E��GW[F�_\�1�\�"�A(��[��]}҇�:��8Iw�1�#��ZƎ"P/1� -}EdS�\�=h����N��8�O�}tl����� ��l��?����޽p�r�	f�����H�3}����'���挐�Q�?=�l
��?�D���f����{dw��Ա���6B�BKt\�4^Eb'�d$ 1avlw$Q��ֲЗ��4ʉ��b X�L�l�d4m=8�iH{�D�*��w��{��@�s�R,���{��g����^w�\;_����$��V?��n�o�}�WI���-$��M��L{֍�eva5FЯ�*fx
�ͨ���b�h|��5V<Qs~`m7�d81	Ll/��u~W� �JK��Nt}�s��1[��5���������)ɦ�bS�$������9"r�xHՋ���R���s5�b��hr|(C)�ۑ��+��������y����-me��/
G�9=����ƍ\&��9�&|_��aT���X0`�,�A�E}yS�F�@�k}���VA���=�2 �[�h��~��#0W�Q�:�Ynp���C�=��F���Zw�1��;�c���S�خ�k��|�G���������p���5���D���&�P߷���x] �_�}uNB�u��U&���:kS�0������I-;c��(�/-ۯVJ,u ӯ]�P�a���ɏ*o�w:�"� p'\}� U�~�Q�ަ�4-�uF�-yQ�p'G�'�Ip��zi�TX�ӿm�;�"c�;	i�H>�BZ-�_5+C�advv$~���d�`���
���!��
��3�Jr�9���_,B���	�f�pCP���^B��>n��~��=j��-���iQ��4&���R�ᲃ1�<2YY�4�)�"]#���b�m&�m��[�%�
X�y�Q���Sͅ(Q����0w�����.eޝ����`�,��yGA���?ja��Ɣ���� �
�̾���)�/ۥ��ۓ�D��#f���!^^b�T���"Ðq��DW�D����Ÿ����n�����N�'
B4�����Y�p�'�#N���]���A���H��}��bEr|3���I�<�� �r7r��`%��W?�Ȫ��w+�f%	ъx�=Y��^�b�%�X���}��	*D/2��`ơ��X���m;�P��JD�'��2���Mϫ��n�4X��c�,"œ�yc?.��g��₟���R�a݋��HEf̀��-S�T>1�$9��7�˾��s����8�؎�:����I��6h�Fs�KJ�y�ag4eFH��;�N�m~(_c�������j�a����U���+��Kﻻ_%G/�snU��t�!��㈑}�|q�>�̎Xg4�z}��"���Xئ� '��Z+��#��/" yM#04��E��䉢12���������ФJ1f�l+c�rM'i��(����}�����Z��Q���JM�ey�=f���{L��B�� �J�+[$��2����	ˉ��bGҤ�G��K��|�� *D����4��0�SY/���➡���I.(��|ȋ<?�z¶�Rx�����`�Ie��{|e
�:p+"y��}�d�a�q���F>�o�F���hH6���k�Q}������7�;�EŁQ Ve �0q�x���b���݄,U�`��0��(��*Q�����zZϻ�>W,�,D���\��y�C�pR��q#��ǅ��y㛔s��y���`��ոo�%_���9(�J@��Uis��灏���R�F�^�����w���)��L�[���'T(�|9�f����>����)8��I�m��︚��-��P�R��H٪�L7�bvl/MCkg�5"�nO���欩�c�T�h�s>�j�>��`a��8P�̍/]��\�ۋ*��~��&ܶ;Ϙ1#�޴:U6�d�j��B,b9�F��,��2��KQ�Afڪ��C1ahSe6��ҸǁR`����1`AzҼ�`8�h���P��ph������k�H_�4�Z$����J�>�Y9yʧ�'.1~r|�I(�U�;���F�y~�;�J�D3@3��`0��컹-*C �����D���o�9K�W��ӣjP�e�;��v�Sw;�Ry��]s@/�N��~�Sɐ����|�f�]��`�t�����Wg!��y���F/ت��/���r,S��{W�ne���b�������5�J�����I 0�s�x~9:R�*����Z�2�gq)���|�� �%�T�C�]ڧ}�X��p��
��G9�m���� �t�>H�U�	�i��6����2d�6��;����fcaX��.�E�IqcӸQ��qȡ5�G���\�%�?����Fz�����Ip�	J)�Ʌn�A���r���ic8���n:����-�BD��v�P�*@X�`��3�}�o��X�F��ƛ~�s����];\pb�<�՜���EB����?����t��6���B���$H��I/�A%�~�E��*����E���*�[(L�􊄆t��6�D�b{¹*7�,��|<�4��Պn�@���z��Mke]FX8��3ǵֆ�.�y�Λ�_K�T�נ:M�����TR-6t�}'�׷В���&�o[�'��bM(j��́J!��xEl�c����gl����^\���*�z�GeӪb���ƽ���� �~�����|ŭѲ�F)�`|
c���h��/�}!v�o��Z�/�������m��|�%��0�\QT�R��������w�w�`zz�0� �G��ZuŃ��"��ulPx��x���ճ�M���]���������7����p��4}T�z��\[R�oo�sB�@�!�&�`�G�O����[9A{s,꫎OȂ��:C@R�* ��
͞Ӂ�}''ʏ�H5K�Y�[����J��Բ$͚��j&9�0hii�ϟS�u��L�2�b3ǵrD'�$�����������۫��"���r�>_�^�Ir<>��G�����^B
�4����m�X�v�3��q�;ml�����eݍ2a������{"í��s�2,9���M�ˋb-������~Ajs�U3D/p��z_�R� �E��)����!3��&�	��\F|&v���:ƃ�����H�����R�ڲ ���l[��7jE����.˸%��!����nr�w�G�>�m��P&E�pZ1�j����l��ZHn�\�⿦ z��dO������j�9�L��P�k?���M|IQ��)zw�8��r���������?yK���PH'Q�����yd�!ݛb ��У�Ӡ���E�6��A@f�y��7�l�E/d�:������y-�09,XĐ��-���ys؆P�g/���@@Ul��y���������7j��5�w�x�D�:�T�6F��IL>�j�!U	��kK�@pUrB2���Jn�|վ5�0�:�XnG21�=:R�g@G�ω{U-�/�}���+�������(�"QR��_Z�
�d9�paf�O����O�SC�z��� ��]1�q���w5B���>R'^�e��{F�o�<���R��{�,�E�����7*�q2��`9)<~�$�M�]k�8���"^HO�đp|�k� �uf�ST̀�[�[R�9ݤ�B�\ �<À`>����KXl�U.j�����T�7,2�^���X���sE"4]�_�+r�^�S��1�L���m�,���"��H,S�6���P����N��l.w1J�o�F��5�o�����e�o�9�k�M,;N��"�^�]�+�����]g�v��=@B(+�w�Ea�Z��,l�ϳ����1Rvd�od����Ű�`#�SJ9���k�����3ͦ3B�̓�T�(�"l$�"%@/}����CvT�8CGC3xQ���}M���C6�(��%�)�0�>|EV�H���=��[����7�Y�Q�3���Q�M,��q;��gM�� t\����7ٷR�Z%�94�d4�g���!�E�̱���W�!}��;<J�[�2 �ڹ�����}(�A8�%�����nm��
kR�@)�ӟ���ʜUY�"�@oL�'��j7�#��J>��E��[����Bl����&�����rvݍt��NT*D������H�>��W|K��T��x���舥'�t6�%�y^��!ː��n��B,"��:������M&�~R`�a8���Š	�q�oۙg>�H���!����׈v_?�KU��Z�c�R����� K���)�����Y>��V��0��ȏDV��#F���yG���
 ���C���m�o��Qw*HʁO���pT�MjY��L��̋I�G�i ?��aHq����?p>����<Ç1�0���VZ�C+F�b��A�X�0�`�<��lP٭�N?)�@:��X;��N���p峩?Z?xy�z�.�7��-��Y��~�_�~�c��!:]�F����x�7y6s�����V�$�MΰFrc�qmЖO��������q�u�]v�P�v?�h�3����� ]�jR�x8r~t�9�!�.�xh�ӡ9��>.^Bo�rD_�Z��P� ��4���xͦ�ث����5�|����(rr�@7J����F�o�R+��:�ÛF�:��GY*pø�-�oP���2�/����.Ϭ)( �\M������8�#͜6��4L"�R�2d(D�ɴ�=)�ӇY����k&V�XY�4��M�2ŗDq�� T�ڧ�KI ���P��Vn6o�4�&�(픻_w pu:���h$�>̎��>̏
B�8=��W `�(�9�*w��J¯J0����)3ILF`�b �t�PV�E��)�!ݮ�2��T� �e��na8��6��h�0.��6�k�S|�������HIPef9����̓[�$�^��4�@_�*/Xxx�6v�`>��-N`��#�-*=/���^y�:B���~��ql�#|{M����-��o�Y���9��u��4�����(}ͩ�h�O�-B��l~0��#	Q�0Vy؀E<5��r�ƨ�D�R���xk�'�,j�-�6@��R]]+$I2���� ��l
Ե��q��.���f�l7�����.f�t�g�+�We	�	������0�\���U�7b1Ƚ��v���j�~.>��RR�6!797���� �2?wF���з�[��aM1����s�Ym��{{�(��=�������̎d��g=I�%H����&S��>L����vZ��V�![F�YM�B)�k�Py�A��;�$��'�Vs���*��OLRGJ�Ad3�����I����%n��K�M�~o�����\7W]���6FG�d��L&�d�<�{�j8&�|O���2ŶI[u/��h=�~^|�'�g_��W����}T?�ЗG�����M��^A ����͡yt���4����(aW��͍��R/Sw�(h�R�F;)�'�@�|ؠ
+�;C	�ֻ��f.y��-t�.���ڦ���^+s��B`�lCB?�����޺��a�����y-<ɞ����8��isu��ˋI����Vj錔U�#N���G~i9���{����Oq����Z������g���%�w�L|on�.C�T5W4��(��m�RI�E�a�NR�z�����kڮ����g4�ie�����\�2+�-�p5����~���mW|��[�;Fx��
VqV���lDr&�TbniU=y��r��z��� O""�(�㩌��҆��rď8��p�H82Ѹ��,^�@cT���E(#ODd7���sl��e�9V��{�|ao\���0ؒa��m��R�>T̉Ŕ�6�XȆ1.pԤ 0����X�}�=6��*,��_I˖ht�!��$jφI�PښM܀�'���m����O�	��EAQ��P�$qp(UB��I��YQ�C2qf)F�:����-�\V`{�^��e�^F��T�8u��D%�c2��w&������q�/���?Ee]�o��V��أA�R���@���!C����m���u��cP��S�^R�а�m�#�sű�_�Ϊ��L�kR�,b��&��V$K���=�l��ڤąV�[#�m���!nF\P��������}0��3z8���>̒�Y`���a4.AL��+����S��pp�z�����(TT���(b�v)l����g+6��Z>���?�p�*���
�k�9�Ex8ԓ��Z6��8E�	�B�i<��u��f�x�p�+�X{��6����]�0�[��˚6̓qK:�S9+!�&�ي=?,��(h~K���豃�o�^�39ɽ��	cd��8g�TbE����O<Yr���Fݕ������`=�V��p(�ݪ$����ŗF-=^����u.x.S`Tt�;�[��g������~�N~'���5<��)O	�x镚���Y����	Y
R�$o
�~>����E���L�!���@H��N����`��[*�H�v�O�\�m�]%�!�@o�����1�l�R)�=?����h��-ka�)�Fw��7_�w���^���m}�/H�5Wux*�j$ ���\�h୾M·9a��!_odį�.�0.��&]�L]�i���G�`h�,p)�>��9ӷ
P�� ��|�6��V˫�ߌ�9s���ዖ��O6�9�@�Ѫ	IF�J�X�u���g��rl���N$�g(k�h����Z�/����=7�MR�\�7�p:Am��N�ƒ!�Q�wh�wzφC�����5�xF/�E�X�Oo�y/�دa�E-���� �Π�2}�
9�A5~�����:T��%��$gTE@M�o�2���M�,��*�/�y4���٧�'SO;��� ��̒m�rb�~�o�d�E2!��`R�t�������]�U��B"�G`x�{�	G,���ڮP�6���@�I2[�-X:�����>��Yp*��L�����z���j�Q���8����).��g�m��|��;�p
��ݹ��9EE�$c�y~-D�3�P��0�8� ��$����)��Љ6�QAI�����#z��/B9��ⱐ?�q�C�E��R��i���1���ᣋT�61�3D^��i�!!�w>����y�bg{����ЂN��w�͘�T���A�3�P���Ot+p��D�?�U�hb�H�	����Ն�urJT͕�^��%�}��ǅ\O�	�A-����s�$��5G�EG^Ke�6ʽGӀ5���f�%|tz+���9���P{n���.��(]��1I��By���SØ���+"�mFAf�S
,@��8߁�*��� qV���,u-ÚK;�	�C���'�"�z�8��h��qէ#���.tJ�j9߼P��TT鸱[W�@)@�:2	Ǖ��TM�6�z�i�D�4.�.�0��1�@�/�z7Jt������q��^H_Eȃ��%I������&�N�35���,YNH�Ưqd�3b�~���T,`�{[�)!���n�v��N��uҏ��P�/`=���;K���J�$�>aD�[�MӷlB��j�@fH)�����hd�f9�6m^�}׈Ѣ"�a�ƶį�W�p�����-G��5y�h��4P2�u4�EܛV;O�[�ZgNM$(�_����x{�n0�[1��{ ��r�\����5����Uћ ����8�C��4��V���0����i{K��7LV�z�QT��4��K�����'-���P%�A����G��O��c|�
����,??	�:�YK��ܱ̄� ��>#~�m?:�_���{O��y_���
%p�^�=h/��͵�:\ z�/Kul9�Z4ήjST7ܠW�rԯ�o)~f�'\�)�g���R0C\�ѵɤQ�O˳򀰍ol)&�����i,�����#6]������7m�T܍�`�`X�!0���'+R��^�T`�_�p��u�a�^t��q��o}��s�-*i�/�CV��
�(�6}~z���-�И��x�;I��"�����6�An��!Di��uI8�eHov/x*�A�c��B'n�VdAj4��l���j����}�ML���- D;e�3�ABC�'��k. VSã��	3�/谥�c����ʑӋ�J��4��O��-����;���ˈ�v_Ѐ^��	��P��}:5�&�ƬU�;-�Y���-��7^Yp{k�T����gv~���c�M}����^��&`}��\�E����.@ ��X�4�M#������HkVdL���N���7�{�G3�mZm�b̼j�Vv��G�\��¯V����@�,rQ�I����m+,ZW.�վ���P<��%s��OBp)��P6y'�#t^�ެ#���lc%�6^���9�\�.�1��t�0�hҁq��6^,{���t��)0�"~��: V�v����}�S��Y��yӰX16�ąG���� �ݯ�:c��v9(�3��Ⱦ���P��yI���H<0pӝ1�v	2ʣTF���Q��BBJ0ࡺ��,&L��	����1�\�s?���T����^W��&\�]�?�M��:�����胒�V��[��gUҴ�{H��	�(�n�8IT��rz23(�2@�eKGN���Y`���|n/�U��+Pb�Q�q�7�򚷅��(\�H^Q�f�̠��o�čtୢ��a42�<1�ؗ;^��M������7��/`�t�T:�u�0�?D� ��[��1����`e�/���f��:T�OǕ�J��.��,2z{fÖ3��{���U�FVe֎�C�_W��\�b��u�%k��3�z|#�7���s	U��S*	�1�<�� v��|��H��z+{������8p4B���j�>}�(�Pq�,�c6d,	��a
5�+g�P�����V&��[�߳jR�9�@�Tq)�Q�N�/�Œ��i}�����-���
�b���fh(=g��ͬr^}���ɭ�ݪ�.�s�
�w�@�E��@���/zP����'��,��1�:�y��y^z���]��I�w�c�4̕��¸;߶oΖL.ϸ������.���+r�kЯ�<�}3�2�<Y��B݌x/r �OQҞ�~����&.�6��ѝ%k]ld�)�)Q-�8�)[���(��෽'�ɯ��06)ﳑM�I�E�2U����ڑ�$/�.� bЊ#�j칁���\�ZAG`p�PjB������W;�Ѱ@&tʛ�z�w�i@H���xI�lH�{�Ch'�:�-�p�X�����(yr��>e��1w�h��rn��B������e<&H��>�����S�L��M!%�i}�T�$����3�tyC��>1bz��䑴�jGwI9C���a�+D�>=�7jnP��B�E��W��g�mK�k,/P���1i�j�8&$�jE����!o�Y�(�w+5�gv��pyh�'5��)P��n�y/�Ѓp�r� '�r�v��e`Wv+�O�eu�lvK�ָ�=kO��p���[f1� o3��c>J��Đ>J�7���hi�Z �V��Kp�`[&��a�� ���2^�f�B.^�I_I�o{�lɹ����us[�Pd6�9��+�z�fgi�;T#	'�9���<[(Ӥc��W�_�rL�_;�w5iS_a{�����w8�-��fk9Pvwd?�<��I��j�-w��6������<�K"�PF���~�a�|����Xs~��*�7n%��Շ�c^���]�,�CƎ�H��T������n�x}��YUs��|�?�f��OOqBCt�
u�dO�82�Tw\p�0�R�<�\[>2hV<8�`��>yD�_����`{<�i����A�k@��}٥�������� �`
�.�y�����.�V@}�~w]{���j`�%�J�r5`e�r��N�b���>Ҷm=!<�k���x��@�pc
�i=����e���![�]\\�}-0��MՏ���*ʩ�l\Z��;�/3�cLA�d���N�%q���9��򏃛R>֒���O��O�g$�U�(�|�-�uy�(WD���;��D���Ka�9�����X)�ڪT�2�?�\^?�J�"���deq�3�ߟ3g#?��,�IC�kl�}I��֧�,�]o�=�۹�_<}S�@TFwO�2��� 9F~��?�^\�OcŪz�;��-��Q� ��i����F�5z�	#���-���*G��7���X�����c:ִ̝<���Z��(���?z(:����ֵ�n2)j��<�.��aE�џ���J�E�������k���:�C:�������{7��1mS`��k%���kz�i7i�`L�����ao�l�پC� �S!�
j�կ�ܓGR�$ia���� v>!zDzjJ`&�x��Q�^S�3��!�=�_Pq3��v��o�,��\�����yY}EBU��rx}�1�fi�if���Q�!>��	ρ�����j_�7�:���ݤ�@�I�5����,s�/���!!(h��a{(�Q2je|�Xii��r�M�w�9�4���m��Ԣ�	��6 �޾�hm��xA���[�f^mi��6F���s^�*��̓��W 4�:+��wi�`�L��$��э��a�<�Y��^Jo�l���Ô�Z�o0��0v�}}���/@��D/�S`_�c�O��"��S�%_�J|��?r%^2J����Rdӻ�Z0Y��q �	���9��Q[·vQ<>�'��]�
����o4��=��p�*�Lp�^hJ��D��~�6"�V���x5'��'&N��j⚡癵�*ª��*�a�S>��;;T�r�R�QhaF�fn����8>��B�����t.q��2<� �1� ��$��N/a���)��x��z<�����攳7&�7�j
B�+ߤ�z*O��!����*�8	��?C�����L�Is-H,�B��s�=[t{������p�;
+gp�Gc�ל^n��\�Y	jD��X
7�D~�J'7Fh$�a����z�0��Ȗ��Y0)��1������g��v{��)�qbf���B��ʯ�7��J��6��e�<��Kd6M������A����Y��ao�����J���@~A���ł��-D�QU�}E�hnbM �E�zf���2;�u��/a/yR���˕�5��&�;���E��F;�dvK��T��K>43A$:��NI��XUXB�����oE�h�k̲��^X>�:4��8#��]��ڱ!�~�jx�����x裂��ko���\���,VAӎ��LP�cCî=A���=��έx����ܼev^�cx�r_t 5z*XD��?Y�rw�n�t�y�!bEq����A�m�i��ŋ�é��2�K���u�n�]cEn!D��ȳ�	��o�>w�AP���B`���L�%?����ӣ�[�*e~D|�\U�[�.��C�3�BB���9f�)&
��/��3E���$�a�
@�K1�a0�Wi��-�-�x8�I9�Xݏiؚ^n�(�7��bs䓭�=��K`�I�vb�D�3�_�m��Cs����!77+j��ܦ��֫�TC(��]y�"�F�L���&��\�*W���T9u��\����Lm�f���s��N����yVoA�b�4�@��i�>��K[_:��"��!j_��uM̫�^�E�l�c&x���M�ⶌ)�Y�[���B�698�y�n�FAyA�@�2��ǐ���G!N����=��fSV�L5���o��G�� 9'���gsU�#C��vHy=G"��	�s���(����n�����)c�e%�;(���ơ���]+�I>:��Rr瑬L�F�Uu�ݮd�ߏ�xi1���k��HQ�iHY/�K�����������������?]�Aՠc4����aGgD����=4���ԟ{5�<�� rEf�g�p������Y8�����w�`�9��0�?E� {n�F����6�7P"5Թ��4I�KAM2��`"���q��M�W}�9�-#ĸ �b�7g%���F{�M�����M����:� ?w����M@bI��jZ�9�D�ױ�܄�6`�����-^֨�_jO��>(�fz�4N�-������xDƢ�j�TH����،~����B��&��8Գm�^�Sx�u�zӨx�(�[��������5�Io����xK�ڟ�/P���=�}Q��d�/\NL�Y.R[��Ռ��Z[���v� ��sv��$Ʀ�uKD�J�ƒ�wUsm,Vi��@�6e����������V �M�&��,W^M���&%ZG�i{p�9EN�]�6�3�v�݆��ĽF�O�;Y&� s�)�:��c���ZN#�=���]���y�7�]����
|��Ȳ��3N��WlI�Wp�!��2NnUI�I���_/����)V������p��'�c::�� W�Djo~OǇ)���������.o���]�����{�ԥc Q��ؕ���X���n����xk��I�,�Ƃ�v����~�`�Б���ѩ��E��t�7Q�HI��?�?�!�}Ho)|�]��/S^�6�@n��VKӳ�`^�画�s�^k4p�� �5,_���邷���w��㶖C�����fخ��������<�|E
_�8��!3�OYW*�5T����!����l�4�]�t��$)��)��T��n�ϓ�C|�<�L+,�*KΞ� sY8�E<a-+��ɚ�+��l�c��hl�Bx� `���v�h��<"9��듸�tݨ<V�wzM຃!����V��]o\s��|�2(˰��G���o�K$���~Ξ����' �Z�Ή��[đ3�AK6˖_8	y9�0zJU�-�mS�4�\FW�<E�P����~[�#����1$R�)��b��0���r�?�̪�/݇�C�߂jǢr2��KX�6W*��6��{�u9Kg��d�-qgE����Lي�0�������{�N,�����<��⁴@���Od�f�p�H��h�^T\���j����T'e�n�Xֈ�F0;��	
[b���/f����2f�/X��hV�qo�R���v��\EՌ�$��[a"�Y*i~ÏV\�ez���Mk��A��r#��g�<F�P.�I�!wSry%-�y��oEJ�`�4ɳ�ۆ�;jJ|�@���7��X��7'}=C�@7�$+9Pǣ�s�]1k�b�!���������k�+��e�(q_��!�Oe��B�ȇ�^ <�[n$��}q�Fp3h���a",�aD�{��y�X'��:�=�/:"*3i[2���{9�ȏ}���πD�֦_Ca@����rǜ��72��f�N6��"�E�n�饜�l��0�֯s/�3�)+�jeý��l������%z���p&���b=��C���z-fT��B³;�w(�� X��In��J�r>�'����7`�����]���l�7���B񞩍*T͑% �#�V���Zb|OA: RX�ր�� ��cL��]��vk�'
S�KG���P��앭j��9mލ`��8�%�#"�k�F�k�;���-��&���9^҂k$|���KQe���%��,n�X��s�>�Vh�#�@)���u�9k��u�_' �ւ5EQ�Ԣ�ö�J<�X��g�z=�g�sY�������ѻ�zu42l	~�N\fk����������=VR��U\�̎#D��Z{}�v�4:7��O�䅌��Df^^�Lh�l�z�L�<� �禱�G�t����K�VfP�12�`4�Q%��3F@ ��9�'����������������n�8"��7����~�2�:]�z`�qM���,�)�Mf��VX*Hƃ��//m�7�HDM�R��뭎urm.�.:
�k��RРmJD�h*�eE���͐n^%;��۴�cNo9� Օ�'����,�`���(%|�DZ;�G)�"�"-�(Y���X�N[�xi_=��F�� ��'VV4a�,��Lg.�lv�\g�}3�5���9�bk��ф)e���*�D|b��������ĸ]��&O��N���Yܯx��5�`T���z���ERx�Eu��؎T��K~�C�cNMH�Q�x[\���:���
�*m<P�V�6�+�3� ��kI�J*���VXhp�ό�gC���cC._G���c��ȩ��:�v��ŧ��F�^V-稖�{�;L�?�L��z�;�0���F.��fӪc�qWG��]TV�\�*�!�S�ϛ�K�3����7�q�w��8�T�=h��(ɥ0M�~�{>cʓ����ȠY���&�o���b���
vO x��h����U�gV�k�5�
S�`dZ��\���N�֭ �z��A����F����ъ ObnJ,�$r+6vn�T�l���"��.��q��W��+��D�~�ż�L�}����U
���s�a��*[�<׫[��j8�)P\ڟGt��/P�)����
�|I��S�J෌}�k���nxq����EoA��:Ej�*���~ϵ1'b�����~���H���4@i�I>-���u��p�
X|}#�o�W	�?��SfE�n�#�����2��@M�UQa��|uf-�8�q"VQ���n+�0/�h������\�=��^W�Jz�}���rV|���~���t���X���O�S���V!m�+BC�K�Ñ9�j�X�5����f�l�'=�q������ :���3�Dԁ|"����݇�{FA	�+cu�d�'�uj�3�Y<.�o�����H��<�#2�.�_��)-����CMw>J��GW7���#4'��t�]\�;@�-��y~�c�l�K}�z�3�s�g.x3G��/��X��KLr`/���[�2d����x�bx�N8i�6m<�(Gf���(�Pm�U�p �đ߅N3�{��@qDhr�崧��@�Iܵ|Z�夨3b�M����4���{0Ђ�^� �ԫ������~��y���^�L���]^*�¡��Cv��QO�
flv@.��7�����L�a�8˓d��,w���s�����F֓۩^n;�_�ʔ�k����фu��J�2��`�/�a�B��b�Wkd �9fz�M<>E� ��b~�S\�d5p9B�׭�b�O��J-^��ѳx?e"�I�V��N�)VJ	'���=���n��d� �):��'	��rb�N��*�0�(jn{��/+�J�R�#�`�lL7(/�	���m�)���/䝍��/��ߏX:R*~w�3����4=�y�p�R����U`h�خ���H�f��O�(j%�?\��2�$bs�7',�~ˁ��!��3Ah��<Q��1yk����6�)�]�f�U��o2��:o�䜮��-��m�&�S,��$l�ws��w�R?��3�`��T_da�&�K�2��-ؾπ�FP:���@�����G9�8�a^6�b�u>h*)N
.X���&���"�¨�r2��:�N߻��ô�r���dg�~���Π�=p�CkO5e%����8�#�~����޴��M�ȶ2j�E�o����߳�pd��nJ_O\=պ�e�|.Se�*���_#�[A3�cSro�$
���z�����8.����$:9��l}�0m}.9��we�� ���w�i���^#tl'����* ��i� �w�s�ɂ��qz�J��eEU�E��������0��m��O�D�{�:E�(?(h@����?0�;iI�a��Ct�	�t�1Q�<i�q"�o�=�5PpM	$���\:���&���:���Xҁ�	�B'-c2}`4���E�h��r-`��w����?�N;b�4��7�24H��h1)�H�����d0��g�}�S)�`y�o~�h5�v�"������G:��)D�נ~R��K�ɾ��� �V�ۯ�<��X�1��Ԗn�D���
�{�~�����K.�J9ɕ{�x�;�|��E����8%l1����Q9��?'�Pp����T�t�,q��l��.hh��a�'s�uv_|䶅�&��5�ƭ����^�U�8��Ŗ7@Dy��FG�`NH�����Q��zLԳ%x��p�4x���ˇm����1R(�@�{�k�B�e�L4��tFeК�J�+/��N�<����R_M��th!yW��ѻ4s��11��DH[�^�<�C�	r�����L[�Y3�P"����8�������5�N�r2�B2�o,�1V��˛&_W��Z�o��{ :2Ȳm�ߘ�q^�ڣX_#h���No΍�E�����7�##� N���6��P�� ���╮Ӄ�{��=� ԍzcF�����bf]$��]�%���4y����Xx�i��z8�Pr���
=|���~�/W�1©52/)|�ۅ&���~���K'ƕ�p�4�.�g@R��D�2*����J�:,�s��>�e��ŗ��f�(䒊V�0N�~{���w�9 �O�������qٷEp�S����r��6;��c>��.т9�e���N�mNEPHy.S����rP`ac���-	��+�k�JC;��kW�/D�w(E�\W�߽��-�yԈ�\P#?s�I���|Mo���,�����;`~t�{{��L�����24�E��{���%�x3�<��VqX�*&���r�@PHL���zs;?���U��`(�/�\�~O���S'#�Ȋ��pǏ�o�ٽ��)T^���o'��hUuQQҦAR�f�7���+���y��մ߭C8	��F;�>{����.px����xV����(�	���~�5J�a�TR�_���$RN�=�)�H��n��N�.�/�٦+ /��|���3ԩ�W�c����8)��L����{(D�܎�<�2A����B���>o�6�����އ���	�5,�HN���,�p��[��w�����=e�	$_�����ń#�ԃ(��*���b��<�(۪��(,��Y��~�6lG��*����x�9t�Pk
���͌K��J�S����IW����7u��t��d�c�� .�A�'���^��!=��UK	����"!���l�_��5pN1�pŨ���k��H��M�� �C�Ӭ�Ud���!��̡U!�jz��־��}i�� ���IAé˅�J��j�.���A�����K�/9��mvE�o+��~���8 �#;g�<�5KVt5�Ě�O��<z��2Θ+��O�E���J�w����6a'�Ж��˖��F1�S12�U�MBXj*��|TPKCp�3�lʻ~-oO�>���-f%�8cy�:F�������!���0}����K�St>�[�T���[�;LƬ�)yB�>ɿ�9��9X#���'F�ӂ>�7���s��]k4��ok�#���~����a�6�'=V��?̱Tr�?l��1�h�d����w
ڮ��Gh9>5ݜE��#���s��
4���w����m�
�Q�aj:=� ��m�����������vYѕ7OQ�#�>ܵe���5�5�y84�p�B�u���Rv8�d�p�ϡm�vN0! �]0�tMgr�!ŷh�6����8���z�,L��>:ػ���۠�\
Q����)��C�d�O͓%Z�[VO��~s�����6����7ŋ�@.�F��7��u���u�-�5�b��/���2K�����R��NW���u`h��.AƇ�FV�s�=|,����@�uA{�!���Ik�8��>$fYof��|�y���7n�'���-�����b(��}���k/�g�}_��gp��O�S�����Z���{��m�"��>{�u��ZH�%��x� ~vn$�4����U�Gj���!�Ee�aoŠ'oߎ�����J1�*�ni��aKx�"I�}u2��ï�;-�W�D���uݹ��0kԆ��_�=K�9�-��6o��L�-%�x�Y;V^����jE���U�R����{a#����'��o�~pY�"Zr)q�~��I(RU�!c�U��l� ,�H�@Mu�<Հ��8������Rp+P�6���t�GXBe�f���ecuIZa[V]{|��U�~���ZA����b �x�}%X|JM�kq$p��A��V�1��]Mz�/1��vO�U�����]��RT^���G��ge�.K��[S���%0_�#���㸵E~A�f�;��X�J��@V��Q>��EP�o��� )͆| ���7�N���W{��Dm�����.A\�{���}L�ɦm)�1�ӧ�m6�W�����W� �e�`O�c�72XI1���H����� �캙'dL���K,�Vc��P̯N����7]T�<��?����ѵo���ֵ�����/����E�-��Y�2��N
a������V��U).���߻!zVZ�t�1��Nd�|}OE�9B���툣w+�>��g���L�1*Ӊ�X7/��c"��Mg�	����V�,�
tWt�ysK�PӾ�ΡR=&��W�)f� �޸B���<�ٴ8m���I�<+����	���X�{zs���M_ȝ$+P�"��Hbὗa�3 �2#T��4VFf0��������z��?��A��~[#�)�W��?��m4:Ӓ�p�?T���j+�E7}�ɘ	,y�1@	yF�>�ߔ�3-�j?#���?��߬Q�U.4�T���N:�N�����W4�go�%�N�ù�X�I7
/�CV�f�o�< �[v�؄v�@���k�kk�>�$GQ�ý�{qR��Bq��Ӡ��� f�<�3��x,ܓ�a!�=�Ua%s��s5��b�dw_��
�@�Ѷ��|��� �QՕ���J[�$���#_�#��z�k@����fptQ,Ik�zf�w#}�}|��Ggx��Y�qO��rJZ����ʌ4`�8�j~���-u���r^���NՌ5��%sHw^M6ʤT�c�g��1v5!���C�aA�� ��]<f�i�c�~��ֆD��^~�s�Ly�ba�]p��ȧS�*�8�w�o|��n[Zm�`W��W������r j̅{\8�/@�G|����s�e;��yvf����?)���&���d��t]�h��P_��ܞ���-�����Je��?�Q�]%��"et-�+	�k��M�a�1\<ypRAbآ������'w�20�g��:
�C	V�� Ǧ�4�>�]���Da��.t9�_��:�`�f��7n ���"_�:��/�o�?��Bv�@A�����$��3H�Dk��wO:��x]��/�׹�n��Q�#���r؃Y�*��u��Ÿ�:��l�Ļ��E�O�[F�aA�����hM��Y[�+�V�U�����\"by$w��0����� �L�	ā���(���	�T�W���Z XT��CQ�=��������P�{�ɂ�d���b��f�����6�X�K�ڦfv��GU�%�Gd<��N�V����	ම�BdV�4��)�8���*r��s��'%�:iӪYݻi��yDT ���/��*~XÍ��}������٫Ѱ��@�e��owv�Έ�Z\�q^$:���.���Q��H�p�>��	��(�F��$��d��68��B�@ii�C�7�C��h��B�icv�׼��[���Dr�s�L���64k�l�����V#4ru�2��P�A�" )e�6��b*3�9nb�$��#�C}�			;�EJ�cC�#̚�=�쾉�T����A#AQ���c�R�֯p���jp&١; Lf�'܅�4P��,���_Xw.
�^�Z��.�\\M�2D���Y�!����H�x���������g3\c!�k��&L���n��Ae��L��ȴQ�,J��;�-�
��B�����:|c�*՛	���!�s'������c��X#�VE*a������0����Ng��D����}.IN��o k���E�C8]Di[M��6$,��Cz]�?U��$	�;+� D���7�n_�DD��X{�%�'�E���G���Z	��
�H-u8�VB_���	�?�����Y��6��ޱc ��lVj�댪��9帕�N� ��˦�����W ��'ނ��omp�hA�q�w�܄n��ޗ�n%���8�^��TG9v���j�a�F
D�=���?�{W8�|����ƛ�I6$�A�����u���1g�#Q�-�<��C2P��PՀ��_��]I�=�s3kO��|Fw�#��{�Jޛ�\���S�����t���%E�$?Sr�T�S:���҅�h��U�l}���歂_>@��F�A��~��v���(�MY7Ų�?d�
&0�.`�y<�-Z���I�%��}4'���>:�Y���דgי��mR��[�r՝ǚj4��p�����>�4�۾1T9k-��
w1�2����Wbݔ�+mDo_�m�I��(mV�-j]�7��l=V-8�l=%��n<Q�d���������ⳍ��� 
[�A���� @p=|W�gF$hC�<k��ǒ�M����7kL�C�-J�W����̾d��U�!`?�1?/أ���H��,g!/_���\�}juJ�Φ�7���%�������Xr Q�m&z��|�4����^VV:,M���$`���Y:?=ϼ�2N��a�� cH�Տ������&P;��=J��i���s{֡�Y�+���d�^*gF�?��tӯL�~'���
sP$��;,��9�(���S�9�;���~���f�MU�kX��L�G�SQ?\��������b,2�R��^�/��nY����'kϽ7�6N|�ݺ���@J@�x&H�d�"�<��b��ꫣ�~-�v,
�C%�:�A�DX�7�Y�w,�q?�/ 	MOd��\�jagC[f��#�"|\TD����z�졁���4՟QOl2(OH�5�S1g
��
�2޼�}�RYR/����n�՘	y�#�c4}30E%G.���U-���- Ą��  ބ��]�\�	��v�������{���aX�Ti��(t�y��C���!�E�U��d�mL�T�վ� T�2��,��5�-�c��ORv�,%�g{�Y�6'�s[��6������܀�.,�R��7W�|�,C�8g6���������Yt�e0p�M��y�2|m'd6� ��#w�Bkg��2���Pjcr�/�|q+�1b+j�mᘪ"74¥����:�Se�ρR+?�5b�z�)�jʋSmJ&+�ox~��[�����-[��bO�je�ɏw�YY��h����`QP3T��)%��L�7q�2�h��z�J���HnFj&<�PN4���(��H%��(9�Wae�!��S�W�=� $IQ��Co%Rf@u�(�A2�/*��stе��k���kW��/��z��<����SN/��*
��Dk���/K�J��������s�����bfg�YI�<ٖ� �[�}%�x��D�e�y���^�J/�HtkJY�p��g�`7r��%(v�eJ���8�Һ�)q����n�����{��XgpX��]w7��6o*{;�E0l�q����(�=X@q*+:nH/۲,+K����_��ޘ)K��E脽�Q6��N��f�D��lwt{�}ݓ �J�y�8��1�����NZ��������A��Vgg���y����=�{,�yក����X�D����pO
đ)�<�n"}��n�:����_���A��2uEl�̹ҭRvh1�� x�֖�oh���vP��	����y4�O�(��(�Н}�G��q;�I�X_8���|��%(�.~/x�4�t�'ѯ�RI�>A�Nσ[��lVi:��_�NO��|�`MU���UD��ͨV@�$�i ��-�R�eFǢRoE�7ػ�$X��:r�)'vOd���t���Þ�=J�-���_aD������Nn���s;Сّ��6.�|uc>}_����FE��m���H�����:�/Hq�<�duFè�4J��Fc3%�(�s�@L6�³�@~�u!k}�Ɇ��Z�qئT��K �����'�ϓ�������V<����.�w�����l"*��r��o�D�1:�T/�驎�n� *� ��,q��>���@�19�����L��3姆7鱻���; �v�F	�<I���*��j��d@��*$
w���A	��ү2�TU�C��#��y��#q/�1[$��@i�M��%��P@�'��R�K��Z������|�,J�4*"�}����Y ���&�
�$![�F7�ß>� 1��a��q�Sً�iIb����G�Aп�%B�w��lzO2��?���OZ&!~�}j[��%�ր��{�E��2L˛���r>��EQ"���+Ws��ɸ^q{i3�T%3~�E����P����->���M�-�o�*��ƭE ���?^-��2��u{��YR�d�U&E���Clo�7��ӌi�6��?�YD̓�#�*����W�<�L3���f ��󫀫���7)�k1CW]6\�Gվ�l�jbs�U��e5�*��7;r��=�rS�=���>)�-�XE�3�(�Y�8Z�a�ȵ��}	�����Z L��z@����#���<��@�+�]���Ԟ&�)�b�:x��t�s���9ήr�<Tkõ����Īc�u����h�Ѥ��}��vboG��ib�O3���4hk{Z�t.]>��GK�G�ī��l�����m2OFW2����c�?nLx��|���VW�&�c��΄�h��� �*��7+]\�qvҹ�� �u$��{6\�tW'� �ܙ�rO��gh�Qh"�|�T�D�F���F�ף�\�kw�eJ>�]��� 9"(�ލ�t�v���0�����5%v�/�`Bjt���oC1��͐?G�K� 0�|(G�!b~�6iz:����'`�']��o����0��c�������iA�9^�B-�̉Nf��:�?�5j[�;S��.��NA�*�0*B�	�i0��g�u�IQU���|�����K����r����7�<F�2m�IӸG %M�7hf�P��S��e͟���u��]ψ�Yy�^&��B}C���������FR�D}rY\ �)"񩃌ߛ(җ%]�U�tL�)���Yr��ǅp��p���%!�I�Ni`z��9�x��N�&0�`�������#��U�`��2��Lbg�������Źl��A=��s�8���E��rP|�
4A]��	�m�V�X��|�D��Hu�W���ނ#�Ȝ6��R&�5�#��='��>�pV�����/�CL�ծ�2��5�>>ڤ�`E�����N����`���v{�e�Ţ"%6w$�ާ���yK�51�e��oae�:M�Y��e�$
�hO�h{��L�	��dȊn�x�)`0������`�2��:����(�C�zD�2 �D�Y���'+����{���c�!����0�[�V�U���������[z��=Y&�a��g�W`'����/2�j���[�D~Isxx��g�ʩ��t�Y��໸�{E�O2��%�ht��܏.��P�[������m���_3���ċ4��떴%	����h�qPW��Ln7����/��������;*������o͘s��=�P
h5���%���m<Y\��l�-3)�^�)���pqC�]��L	B�3�d?���d!�U�a�h�yZ�ƲE�M[֢.��}/�fo�cN�U�����U�������D9l�]�`�#���7�዆ᢀ��=�I�q'���M�]Qo �)j�����\ku�yYSD���?ռ��z	�oz-�4��eV���G(�WP�&RΜO���!��(Ha��,Ż�w�e�����ߟ��j@	�L�6�ɔ`��#�����V�`�1c�Q��(���,��3�v6_%+����bҌT�S�-
�o���ܯ��;]�Vβ�"�J�2Z
b�)�X�o/���C�D�x��0_��mw�1d"f!](N�-`ERK�}�/g������+e"��-"F�@��BL�U.{��"�48��bYH�{f�Z�������n�o������f�FIN"�`�H̏c�}n�6�0��i�m�\J�VAm�D�mτP��f��hҕ���ϯ�����j��,y�c	�\�^�x�Ct�-�����r9�k�t��+�}19���po\=�T�Ȱ�t������Nn<xm�oe
�y��c
�cV����?v��O�#	�݁~�U��I&��ק��Ql0���ΤnnzЅq>\�8�W�5_4�eנ��qCR~{<,.FL2tЊ�G��h���0���^}�'�&�u2�)�(%ʞ�''��zft*~��74o����j6���=���=J��3��._��s=?���FYU~�F,J��DC`H�?Pi�L���"C�_&���w�K�=0�Q��_~N������5������_>ܠ�����K�豯d��C�m�pe�]�d�:�+����H��N��	Ѫ�;�jg0 ��8���3gG&)�g� {�L���O�)�*���y�()ԞRը2S���i��'��ܲ�'s���n�e���D��F���Bx�����y���Lk�ߚr<��説z�m8RBÑ�����uӭ�C�R��[�zf�5`�&"-��2�{Bw��*[{�����ے�!�U��"��2�3�>O�ܪ��G,���Y��*^�0=���H��� n*V<���4�iXi%������IX`ѷ5�İ	P�ϯz�,�+��}�Yq8%@�\w	:\�մrg�R_b�}�GJ�Nt�Rj����K��u��6k`?ߊ�搇,EU��F�o�B��x�Xk*$�A���$e�ʨlv����_mw3_������Ō�O�$Y��l��6���܁�!^�N˹B�󽁶%B����Ed�Y�i���qv=�g �/��tٰ`�m�n�h�ܒ$�����T���NzSб�!�y�r5��逇�}ߎ���O�D�n�8#�Pk!Q�O�"�g�;u��5�p��Oo�`Xy-ϩ7a����i���FJ�(1-7:�H�F5����rH���Tu��{���
(�Y0��&�νi�&��[I��x���:�8���0���ȱ��)��\��,�,�։��$0ޒ!%��z�Ӷ���\��@�(�[rJiV'm��؎v5%.a�ʊ�H��۱�sȴ�(Q!R��u^�@Nm��_��3��[�"xS���t�X�HP�H0�d�Ɗ���>�"!��1�h:F�>!f0K����y�&׼���}��:�l#ˡ��4@��5W�v�q���0LP:�����F^�_P�B-���4���c����h�y�?���O�%���B#�u��Ie�;�]�9��6_�?��Q��.�wY��A��l�"�CFrS6?��E_��.}&%�"�v0F<4�u**���zo˚?�����+��=�
�ERNʝzKo����.���TT���_#?��.��R���s����r0��.�.	[^:E͔A�t ^�p���T�9�k6����v�;G�[x���$�Io��!20�<D���k�J�uBa�Y�3�Py*����U�=����I}0��L�8L�H�$��`E�D���u�.�_8kڤ�/������C��Y����3yFN��LƊC�M�9��xe�K�9�ߏ���3���&3W�%\��X �ِ�� �ʹ�p^��kr{��.yZvEt#e�h���f;�������sd�pS��yF��	n�U��ཁ�i�x��%�Ȝ�2���6��N,��8Y�;��2��+��o!;p�sN���ˁ�m���L��
+L[����Q,������mi�����<�͑߱��IK��=��k��:=��#n��?_���߇�K[J+�ՀQ�d2R�M�C�_������I/�j5�x�I"��F� x|7C���)'����?�&ӒS�U���uo�2����ӷq�0G����Ai.���;F�����Q���to�w��0�&�O��o#�� "G�� ���kRvd
eͯ>���h�y%N<	����a�2�qcp-�|Rڿ�w�����zW�����w���>g/d#�#A�BG�FdX3����|uf(3�bk�U&�&�4�m�����]�TJv�M�͊z��,P�Q;��� ����0��[�*j���6�4��p��Jʍ����3(M���{��p��\N����?�?�SO>��'a��ޔ�JZ�)j΄�GC�mN�
�Xr�!�r\"	9�3?u*1�Wlm*;����	}hJ������T�����_9Jp5&���9 �-ǭ�b@ 	K��}^e?�������w�C�����C�o^��h!��E7�#�	$�o{N�yڂ^A���X�i�~��$��ry�d��<X!����q��JvB��vp���-Ke�4�qd��_�rI{��%��.��~l�=\v�=�l�(�ĐS��A�E��J�7s�>͂���G� ��B�87�>�EE�[?�u�l#���a7)�����q�&Z��T/ۧn���_͂��U[q�1��&�K����J/�N����9o�g�m5�,_|��pIz��sU�{�0u,!��7v%?�
�q
�D����Ս:�}
v����NDu�RgN�������Y�.�a�a�H���[ k��C��~��[�b6��k�U��h����'�Q��z�h.���N�p�t�J�O��}�E�:`���� 9��1���?�'�qr�= 3�����g;��WY*����=1.���K����d-K|�?�����{PkH����g�	�`� ��d�x��_�q*�#Qp/�@�
�7��4�+\����C��H[9��5�<Ol5��h���3����蟫C�t3��Q�':�X����6N�����Ɛ����;�e��V����@�-�Ɨ�}�"q�Z?������7y�=�u�5��e�A�a��L��?����ge�sp��H�oZ2^�w�=�'�-��O��I�����^������h�;BJ���T�ҕW���\إ����b��|�sT�ޣ�g�����Ki��IMn�p0�U|+�nOn9y�(��'�\�kSA0E�� ��)��A�I�W8K��RvZ�c4�$�'C�VC���j)���?���5|Ke�'�]�0���v��H����(�{H�;y��G�R�Ї��*t*�}Qg����0¶㑎�h��R�˄���~	N��|�g04pR��޷��_�߷,�QR�BX��;AE��c�_����>����l��7���}*p_�1��8ڜx'��{&��4$�#�EA/�]��vM`0�Lf��ۯC�|$�s��<�z��b�O����WM�:yO�ԧs�Ä\F�'VҘ`����AP˜��K�E�%frߛ�07Z��DwŚ���+j�J�����6�V�����f��,�n����X�8p�6�%6i��Bzg�L��ʙ��LP��ƽ��J�[���V$�	H���o;����@@O
���T�2�`|��٣|��s�h���Gb�7�i)�N�c0��@�9�T�^�?[����>��Z�or&O�iY�\ �3���\��$0	�f��8+�����I�)�3d8�.�q�IkKZ��Kz����O�L>�������;��%/�I@��F$YL�Պ�eW����s�f"�/ŽѨ)��Je��q��ɂ[��V�wMR��b��j/6b!�x�J
z`S��Ҏ����B�ѡ���(�Fd��DaԿ�yq�P�l������t�8���f��D��o�d("8(VM��
 "��M�6k�W��B�	b��&�(ƃ��rڵ��&+c���z���W�æ�7�����ň���+E8������f0*|�!��Q��O:��zbι�Ȁ~ߋ�jQs 7�
�Zvǁ��F�wR4F�@q~�4�!�ߴ�ٻο��f�nYzw�|;�J��G�/k�ȝ����yQ���"uX}4�S�|��p	��=�"�7��;;_5��bH{N���g�ߢ�����K�PW��L��h!�@
�Mq��!�F�Ĕ�5�����B��aD��V�#BJs��q�W�N�r����)�?6��
`�	i6�
{��T)V���;�ۈӹ���]!�̺����^E?�quuPah�(��O|jr�*��i,�xx$�Y%��9ඞ�SJ�i�'��!�Bԓ�������.D~��nJHV�׭�9T��Z������3��.�3y�L��	Ƚ��	��M1I�.ނ ��J�U����F�`!δ������miY��/��ļ_�lZ-@2���O.fp�:��]E:jv~���?|{WG�糍�^�����R%
8!X&�D�Eb��2�N>8�����R�;w^��������������`����b�9p�ڽ?9Hf�Li�RaF��F�����	3uzF�	Tc��]o� W.g��ō��(���Z�BЩ�,��M�l">�7ߧXH~������WO�2�K߭rР~9�nhW�/��9$ݫw�}��Uz)_ꖕ�UR��T��b ��͘�Fo��yo�1�;?�#o�k���,�d��^.Ɖo��G{+�m�S�l�u+񀥠��j��G��<�U(S������T�O-Y�X�".Y�6D�t!����� ho7�; 6eσ��[V<�iubG ��������%�
�Q�v�J1cٳn�<J���=Hb��t��\�7ѨN<*'���{�*���m�����%��;1SW�崔ڪ��e.�d�<�����/���,�1
�,ךޡ���ѩ-��g����3��ˉ����Ի&0_#h*(�lq�or��	G�$[|�L8��i�˹p�ͧY����TS�&ʆ����^������1��� &#xg�\�74�a%�m��ӱ�X��ɪN�����=ع~w���~������y-��3�TmQFI=�Bpp�?EP�x���}7ei}?R�F mqǪ�;>��-�7>Q<�T0Ȩ�3�'��\"Q�ޑ�뱦,0��«��([!�p��L��X?�j_C9t���i<�"�k�fb|�T���2�C�[��g;�bYCeG���
1lH��e	m��D*�~��#B�L>Z<���i�A�-�#���sT?Y2J$7h��^2�����;�,;�5�%�e����X �`�Mc��E�7�;���᧼�I�T������p+F�$�'�&�Y�64}E2X����4%�����'�\̀��0Ԩ���"�2�G�ֶP)�G���#�5Xi:$0�n�C�JZ�����6��^c6y��R�U���l�ji��F%ȥAKqM����⨓��E�C/6�%�G;�u�%1��R,�a�U�%5��E:6����1����E$�<[A]sU��>���}}#����)^�F0#yU�G�w�X����KQ���{�;k�Jn�q�\Z&n6\,jb���졼�m�n����TN�ov��y�Fܼ�k7�uP#iʌ9h�.v��9rz��7�98*�D�+�s-��|i���.e�+�+�2{�Д�%YI`azi��ǩ�"��2lI�@i��7mD>ㄏ���yK��A���)s���RM�=`9�܏��x��X͎ q��X�Ƶi�7�OU�
���4k}�|[/�.&�@]n��m�:�q�1*� Rɨ����E�7�
����Q\�ˀ&4����<,�l���=�G6�ԮFr�$�Vg���p���j2�@?�E��Vq�_{T��-	�*�$�?^4}4X�A�;�Д�I2�7V��q��WtB�4�~����WL,�z�([���:��+�ӱ�.�;J�h������i�Y��F/����	R���G�@~Eu�e6��Ο����h��xI����C�%����?#�]�����JA��pD�`6�����=[�pU�XH<u!h젙���$�#����f���lI�Qtw�oqO&���U��کv�+��,�;�·��0����mZt���M�,e�,�K��\�ǎ �a���lr�r>JDa߅ٜ�Av��P�X{����X�5�#`���b��B�,�P:9���O��kpO��l�
���&K������mƻg�m�E��FbH�YEfv#�~���xHI��
� ���2���"��z10��h���0�xeCɰ^�Jp-%�v6��>��j�5i�o�c_����
ϝ�G�0�Ƹ2�� ��Q_���@d������D�G�$�?SD��R1�[�U5�b0���8.��/����0�E�?�l��l:��oh�)�	�2�����E$pe�n����D�G�m�%X*�K�?����C�^���Le����D$
$�;��eV�A�Y`�kO-������������d2r��$�T���Y�����hq�_kr�t��K/�K''�P)t���}5Q�SQc��[<4�@�[�P�#�}���@��hy�b� �x�!��*���K�`�5<}+P�S�m(HR��kT6,��a|k�.1�����r�V�F?�'r�~7Ѐ�=|�:oR���&��.H��:����a���,���S��Ȝ����鈋GD��F�8�׻��b���'�H7�G�ҟ�`X���Ģ���,ۉ8�V�LA��E�N}�$��Uqw���\�Ý��1F`�fc���R$|m~P���h��M�#>�8���ˉ�V;kYIs;�x��������K0YҶl��z�2d����7�v$�%f��de���7DH/�� �X�Q�f��ED���d��W+��%��弍����?�[۹��s�1�(G�P�6늂����\�[
�\[;��!3|T[$ͬ!ne^�U���E,�k�3��r��O~���_���#W�35�#�3|��Q��ji����f�����r�zJ�S��лHPK6�]���Eu�8��P�v�C��s~EhjcNW�K�	�O��|xUZJM4�hؑM59׏|�C�Y"s��K�وF^�*��Qn< �3���<�`�����ؤ0��J?]�L�&�(��	�3Lû�
T���e��D2I���YW��)w����E��4d*�Q߃t��/��
���Ź5[�G�����YE9�}�
0�X85["�����x���Z�3� ԟ��y6"�ߟ*W�ju�Vi m˥c�1a���8P�Ǘ��5��7t�w��E�5R�����:8���C���6+*9^AL�a��ZP��f�R���_lw�a�K�q�Ҍb<'L��G�Mɛ(�!Z2츻4�^��m��\t�7�{��������7��j{Ni�/ҩ��=W��4�X�.��)�i�N�e`�@iL'hԴL�5�����_�$���;��n6C�� OQ �\i/ZO�$W��W��`3�z0_j��촒��i�\ۢ�_�К'�Hx������-��ϧ���]�］�����!��z�������{���d�ꩶ�� ���`�����E�nh�L{	���$�)���+�U>�uP
[�
+]�R��L����7�|�'�L냶](g��<��q�`��^p+�n�p�[�&�J�����q\	 �Pָ�)����Ě�^��'�ȶ5U�@� 3 ͆3�{Q�I��}y�!�G+�>���A���MD�vx���X|ϙVn��g�q�� ��񆩶�ƀރ� 1F�\s�c@^�m>���`���J�2�(���Jt]�6q��І6��+��>Z�\����h��|��V����LX�����g�ʕw�T�zJ�q0Yd��ll�Ȝnt�fs�Z�5g%����PU���I�[ Z�Kڶ.�-�k8�bY4sa*` hE���;���~�=��&�-���S���)�c�jA�� ��ZY*|q�v���Z���#���q}�)_��k�8`Jw5��F2No��j S�p��;��
Is�l��E��΀i�C͒ղ��d0�2�B�����3E x$F�k�Һ��Z��=�l5F�]��3���X�ў{�#��y*��d�]�Z:�E*��H�4<�h�4�����܃%�g���ˡ[�YxQ[k}S���f�t ����)�a!�S5�7�4��8R�B��v���[��#<�&�	2(3O��dkp`����$|��%�|����o�����U��f<e)��j(o��;!#��q�Z0��%�/�u�8�a�{	D1���; ����,'9<V�`���Q8���wH�`�� Tݶ�ߎM���VG��r@_./MU�8��ܐ���	���vF҇]���8x��s�!�yu���~H3�GK�C�?$���G@ҳQx�'�~"��u�$��͞���N�DN�+-�Fgd���R_��#ݪ~�Ŋ+bUYDS��"�{�G>:1f���-d%�IB�f�v*.� ����Ըr�^ɳ�S2�.�����/|M�"[�Ƒ��
����znd
�c���H�L>� �yY��&Qf�9�Tk'��	8]A`^�@Զ݂h��ږ��u�c#�/�ʨ|˩g���������4y�1�7�o�g^&�~�9�)ǕZ�7׍�sa�?��	b}Эj��*�*��p˃#�NϺ��ǻ���s����qp�1�P��#U��*�tFTw��'�U���DO��Npy+w�B�L�A,XUH� ? ɕ���Wq�ڊ�<WΡ^��݄�ۼ�s}PC�'xg��d
�@2;H=�������W%�R�P'!���T�	�$���d	�͌9�f�/p'�"���D�KdS=�g����yV�Z"�v�A����	�*eۺ�LѦ�;��`ҁ�8f��ogLr_���"��u��`��X��&�z�`���w�`F�t{=5����V�ari�z����
���ʫz�aW]:�a�˛&�X��A|��`s���,����%�l��b����آ��@*"��zie���L�!�S,�<��r"��X[! ~<�^�e�UE���z/;���_��X|�r(]���s"}Y�%Ɔ�2J�ڏ�㵔���"C�펙{�S�\�ÞϽ��I[��n�%8" �Oe�U�b��h<�piO�~�B�]Hr�7﹧'��E.��z2�>˥�Vև�����׿�c#��!�?�?A���R!vk�/5��1���l��Y��+����:�5� �B�lk��al,ص�S�de �5Ȓ]���m� V2U1&K�`Ф�f���U��� ��Hq�_F��ea��e�=�%�
sޝ��*�"0���7���M
��dZ��M(�	��Rr�ۖ�lOiSAlM_=s/����gd�O��U_�M�^)muH���<����F��ޅi�^{ �g�\g�?�S����	k���9;��L�%�6�8P��>ʫ�q{��w,Q��O����/�����G�����z1s��z<����w�ݬi���{��#I��x;�����e4�jre����e�TR�Yt��0�1�q�9]��L��lN���</e�^sJ�/�d� Ϗ���X��ٿ5mT]Vd�^B��M�||����hpGOd���쓛��Ljx(��L����c5�����)R	ޙ�=k��u����'�T���PF�w������r:�9�z�y��̸Ux�6�������?�A��H��bJ� �a����6*�x�,.S�:c[l��l��s������'G� � �G������p�4;f������U�`(T{�Z��:(v�c��MZ)!	A	�jՄ��ȅ��=z��QQ�mx~\��T���o�B{@�Ɩl�L+ d�Y#���^)�s����<� �hl!�9t�|I�vL��[���&3-P��,I0(ig�z�����S�u՜Z%u�_�Fo�J��9�\ͱ/#0K�BI� ���C����H���~����4T����}7�+�[��#��x1��secJC2�&��P�e�	*	i
hd?�/k��e��L1z5�v����7i������^W�i�O.J�������RHI�{c�SI�{�e���H���p?���x!(�|���K�?�+��:�l0z��H�D��&#������5���=vFs�^o!(���ڳ)l6��<	������g���龱��I"���	5s��z�� �\���)��JX6�W�94�+�2�ª3'c/��(�p�s/F^�X��"�w��h��p�=�s���ƻ�JJ�/��ʺ.H.�"2lll�cG�zj������zp'K���z��P�3�s: S޹l�}C$[�H1s�?���b�Uq�I�7{7W	->w���Vu=Q�t�d7�.�L�{�5]*�4o���aݥ��,���b���WW����G����4�\�#�.r��ؗBU��Q�0*�߲�z�&�:ߓN�*��A��[��w��'(�#�$�z&B�F\���ey@:�����hO07ƅ���dl �dE�hʇ�q�p'&�9i����R2&Ӳ��z+;���7f<r"c<��a������e��P(�o��_h��� Ƨ��,+�8�"�&�׭)�����,ֳ��W��x�=�t�0K���A:�w�Ɇ�&~�>�D�1��y�uiɝz�䙨�k�/���F�"�0���
�,��e�d��H4���?��٪���4lU��í�(ͪ����	���;�@�9vC�^vF�)����@]��ȗwBXWp�kIS�~@�=�xg	�]a 4�@�g\!)a)�j�8��Ge�Ēi��.δ�Ī�t�����7�n{/߻Eڸ�ב�)ԑ-��8q�^�jg���1ZA_���Imf�M�8�ס$�I8�E��C�c0��>�n�{���e���jߡ��Q�2��I|t��?z==!TV�Ƚ�d��K��6s[c;���~�[���Q�{X��p���*�P������j�[\������H�n�g�^|G���ڡ\�1�y����Xj���ם�#����b^d������<��i�q�mO�Ԓ��Kᘿ��l���e�!D�9})/f�!��0̻s�!�[��S�A�(�~����O�х��*<]
���S!�b����]-(�FF�I�f9��pq�SYV��]-�&t�ǆ�02 ��P��Sc�{L?O�Nj�J���.�g�an��5��,1E.4ռ�·:�VH}�<�12U{zs7tqc��ԒrY��4���n�f.�#�JPq�|ֺ�52{$;��ہ:�|_N� ��d(�ύ�6�s���z�4��׳��d;�)��3)1C7C[Ut_[��3��lT}��
��SC��苃�� ���E{��#��� ��O�!��U�&��d��1��Z2���$�{�x_�W�x�� +��g:vR�?���5����%�џ�j�N� �d��x�mtt���bYR���>�9 ��}�,���i�oZ�֘��, *w��d(C޼�S3�6�U�i�ͣ2�)"<��^��6��%p�!б�a�ZS�l�nw �8\:��W�t�H��!:};	��.8�a�R����+=l~�_��w����I���),Ҿ'�	�O�	s��/u��4�Z���V��>,�O!�P%���F���E�������6�&���I���4�����0������h�/�@%m�+��n$b�
,�9�B��T��kz��2�u�ޙ���/ �0�OP{�I��NȎ�:UD�A5V$rI�J2�u%��GR�Z+2ǀc�@�����
�k{~w�:�&��}�P=�,q$= ;���>�'�8	{���D�X2���Kw���z�I��aW���IyV�����$�Wh��ᮽQqlH�oZR� g;D~z5U@�)v_hV��Et568�~O�
Ǔ�s�^����h}�3}�s^�h[Ue�@!�b�����1��{�O�E	q�: ��$wi���{wf�{D�o�ԵTt6럙��6�u?���){���:������gx+���rۏ�Юf�Ѵs�*i�T=+��&�ز�=�;���-?��k�[7R|V���>�E�<x�5V�ߌ��#����+�o�v����i[0U��QM�����W�s� ��Y�����4zpޑ�MS.����i|�ܨ��"�k�p�/�nm�D�Y"��7���DѢ��|��Qv���� w�S����ۣ�&���.�P�
�Z~���0�=<�U;�5r�R��q@�HiX��W����<v���@J�@�ǹ@P��ī2$��h�谷Zp�Y��'`\�>RZE��lAZG�"�NwhM��,���:q��%��24/ٻP�ZP���F6"L�j�<g�m�`B�&�����U�2��3���K6|��~]����@��(�� Li�����ĳƩ����T�:���̺P4f� i5����,q�z�!0�z����zz��u^��e��N_�܄?���.: G2�9�uA2?�{OLL<��l(@?Q����kb\I��"�y҈�j���ԆU�{���R>��j�ݎ?]كp���9VAq�r)�+Z꫋z�fG����D���"b�����@�S
����a-�G[�?c����)��fe��yq�xLnkv�(�z�&�v	����n��c
��b��\Э�OT�#s��EF��a�S)<X�h=.���m �/���W�4�?�m����\]%�s,0�˘����,�	}eT�gO.�*�r8O��<7 ��oM[I��H�s�(R"�������f���}b���<*��:��������;�
9=�=©u�<����!����)#����)hp�&��h��k���k�A�d`�\�\K�1���gj���D���!L��b,�c�.g����<�3��h~��<7N�;p�m"	T��X1����"\r�M���{�v�g����j� |�ذ�n%p�S$>��u�n������h�<5I�I�fB�����"�A�&C���̟/3c!d%��x"��}g��*��q�0�6�2��G�C1:�� �ܨW���RuB�*���n�ϻ����pb�>5F!��'��D
l,��,�ɛ��	�v��	��S���l^*B����c������A(v��`�ȣ!�t��NA�����ET�`�K��n�9�c��c0�"�Yz�_��zn$��`(�9��j����v��:����3ZIW���55�5`����1�r��h��;�)��F�R�����U^z���tUoG�X2���g�W�¤6�ʭ�_7��4�rI,����`��Uky�ˋ-�-[�؎�؞�C	0:ҾAT5B��[H����	t����'Ďo2��^⌮<{��.�;�6�Uq��>��)�b�V��4u�
q����iO�^�m�#�)��'6GXU`���G��+.�>��>vÚN(��4�u��Ǌ���,�&��2��S��b!�茨A*�OI&�����b�|�p�C�5�уL�f*�ة���������a6b��������UP.��vhyۥ)�
iڎG��æ?��-�x��W����SY�OF˝�����LՂk���L�������K{;��B�u�{)� 3��R��1��Z�,E.��?�FI⿤�=ZZ(�� �j���T%���}�����⻨��xS��t�ᨼm�9B�,E�� ��4�6�d��C�mg����i,��B�jA�r��o|��'P>&��7
]2#;0��s:z3����7�V!��N^׬Q�VU���|��ʦ+�֘��lB0&5���ϑ�ς�%5�%����C����#�M�7��Z������]�p� >�Z�~\��ф�^Qr��S���@���^κ-���F�vA��v1�,�7Ow\����z���O.��;iu�\��O:���<9���t}�b�ف>8��������'��Hk��3�[�a��e혥�r0�
v��'�D���,bc\��x��!�|��$6��n���Ã)�-�_������*��U�c�UjҚ,�KvQ<p��8o�~�*L�G�-��	����Q��v<�,i�j��/mD��aݪ9(��%"�~���8�����d��H�$zPx�6Ns���%o<6�F�}n�Y�HsM�N�ƨ����w���9�O�uë �O�l_�^څ+3j΅�%c��(�����Z�T:71
"��g�W���,:6hak~Z�������bC�V��*��s�H���5��\ð�d��8�����(~�]WލA�"��`LR���~��wM���n�V{F3ؘJ������Bi�e4�"�C���c�_�E�V�����$D`�cgCR�āL� ��Z�{U?W:3��@��T���SLg���(��eU(��H�:�}0i�uOw�Y���4�O�ۋʉ���$r6���兑��n�;d��-����fiS-4NH��Mt�%�G��Y�VL�c�d_���+���N}\�o�3V(F����	.p����z�˵�B0�����>��N�����J���0--m�vϮ)l�i�	Ȥx
�$�[��!����t��Yǌʆ7�a�u��}ë�_��,J�i��g��ξ�vt,L&��@�߻��>�=�-�y�"�q=U�k��XZ����	n�nx�4J����±�nöl��yMn�
 R
=�rǾ�h\5���:��dh��&TN�=s.W��ݷRa=(�ZO6D>�!�J9�}<�5]ʕ|f�!��W型.���v8v�{cͫ�B��u��׾�R|3�����Z�@�ٻBI�ly�7J)��)� �'TR�u����M�lf$�SH2HW �D��T.�m�|=E>�N���IL����"L9I�͟j]#��[_V�¦��d�U������C��S��"�	z�����H>���F,��h 7'2W�<F�����8�}�<��l���n�$u�Fv7��L�9�X�q��n����(�C�Ok�� ��밆��(&�Aߩw�,�u��i�z����t�̎�tÑ�"��~����(�����r��*`Nmc���d���|A.&���o���|{�o�_��T�C�y��.2��̷��Ý���F��F-����Ƚ=����ˑ���_� q!Y���6�DQ�zd>��I$r�z�Z���=? �Э�8^����L�5���S���QX�s�u���Zj��,^c���e�?�C�@��@Uc�x8N��W<;�o���ܕ�]��a*�~ci��YT��V����b)N����g�xq!�����-n�W�����9�!�f<cJ�����&��`��wZw��;��sJ/��:�qERkm���ǀE�_I@�)4�0�����iH�4�c@׻�P	'V7m�렯�.3�%����y���A� �Z���S���&אa1�9���m �N"�`5B�	h�!�ڈ��-w���[�Z�t�I���P��:b�q����c�}�°:���5�j��$�3X�Ն�9�&_}'�Z$���:j�˘�(5��KD��8�n��0����nMw?dz#Z� ��W!*����=��ZD7" &m�X�;a�䪽�����r̆c��-�%Yo>.q&�mK������W�\�6.��͠�&��>TL��6W�s�87bI��6|����6����,�t�Ḫ̠e]���P�b����i�~?����u������LA�����ͭY��&���Z�ɗy����珨�>�Ѣ
N�	�)��΍5� #	!R�E/u-sj�r5P��|<�D{e��^��Q3���������U$���Ƴv1���b����C��'�q7�:���ڥ�|'kO��و�&��*����[ �;����%� _�1)��d[�@k�ȅ�����>'�z�3�*�?\�o/G��ʼ��:��$q�ze"R�;Th���!גa��.�s�٦8C�q䌌Y���]2zeݩ���G��Y p�T:n_	_�7(^���ϧd�̺\���j��65ؓf���79&����{���$���u�z�+#��SD�x��Po��	�hk�6Pu����:&B�ތC"}H���Ɖ}�yKt�x|t��&l��Ys���Ɂ�y#׾G�a	u>��r�p rm\��u��%wd��#�C��.�^%�X�:����^ַ�dk�Ξgs�EA�m'��)4�O�_���5����y��[j0imB��k�6N���0�� �n@$�Q �im�82���N���:HQ�6�QG�9�N��$!;Clu�Qo�Mfw'e?p7P}E.>2Zى�Y�r|��>J�&��K�F��*��g�ǴY������x_�s�ﺮ�_$G�s��~Kk���\]_y�\��L��薒�.� N5�Bb�1�8s�[�~�崄��A����so�m{�E�����] C���Riۿ��%�`%r,5��p�����GJ�z�V�S����~�ߍ�~k��-����rtE���)�1Q��#O�^[TY��"]�!-QF��Q����Y3�;�cF�ƅ��b�Q��R1�%��:;CS�n	ù�38�DB/߂��`�ӏ{�����)%�W�f�n�r�6�	v1 ���P�$���s|w� ����$�h��>��|Nت�;�8/��z���iĔk�9t�7Rf�4�B_�����-[*��ի�_�-e~��;��q_��<�.hʓZ#����Ø������<M��̰01��n�g���G���ͥK���:�ʺ���l��TFi���Fb釜Yi���yד�����܏w��l�	�A�G�k%�Y����a6�W(�[1�_L�_i�-n����C��pZQ�NQw��s�]��
��qE1�޳yy�_'9w��L�	>?��u�,J�����xI%����!h��UU=db��p������}p�ތ�\��;�H��23J�ȥ� ��C�@ø��Z3��p����F��7N׫$�t+��I�Ek�{2��p".,f�꜠�5�|�6 `��
j�בe�p�'V��v�ȟb�J?�)sc���<E�@�/� @&�<B�� j�/�8�ߺ���k���;��]^!K��M�l>��G9N`��?UZ
��ݲ+,socz�n/�_��NY;M%�]�l4{�ϸ"�� Yϭ�������As%����?W�3���VN�����ؕ[�e�k���z@�.�	'݈
z�	�+t�˘���JAuU�|p����"�3�-[�!�|¦��	�ĩSo�ɯE[$N5�9x9��o_	���Y`,�����(�
|���;a:��L��T"�Hy=s��2�]�'� ��
>���E�Y1�)�a(!���d"y�6�pj���F�9�����D�-���� u�\�����c����riqc��m71�����sբGbԮ̱�����
c����I���ϼ��Ŝ3fp�Ǔ����;��������� �f��ZIXbo4���7ښ�}[�8����;��+�j��W��kdɒ���B�Na����_�M�c�3�N
���צk�fN��O�h,t��N�<��	���N�o�]�@�ըD�Kk7���Z�&��u kg�{�
���Ոumj�\��k���i���-T2S����0�&:2�@$56�2��������}���&Z@�����8>�R�{����M�Ʋb�U ��;uV���w�+��	����+���s��+��P̈́�/�Mf�@^:Y���T��|����y�J5V�c�2.-���֪��0����m��9mH�F WK��N���jZ��u��*m��kb��-�V�]9��z�Y�<c�2����D�V��O蟸���Z��Sx|�d���T��Y{���i�g��h\�H!��/�g��B���
�3�az!��1r�c��O��8f;b���(E��!��j7��Ǣ��Ѩ�~�l�(*݇Ӽ�֛s��h�u���B2H�� g��˟e7j����{\'��������UO�#{������%�oGިy(�%���/��$�D��1^ ^\��H%ZGb�}�!f����|_��b��5����&���MI��a�L���O���lc@�5 2K�H�Ao�`ŉ��X�(?��p*v�c�y%��ɑ�a?G�3����R��_H+M�l��"5���R?�ݷj��j���8��N��T&�xyV�α�ޠ�+7�j<����ci	�Z��
�.q����H�"�p2X�C�	��t��#���]0��;X�p��<%��� �y\�t8ITB�425׎�����sbK-�c�cc
h�9�=�e�N4]�Њ8�I
~����ׅj: ���L���Ihk4��4eB����dN�1���nL��~+
�T~2�7��0�?� �ӄX���W�]�7D%45fO����L?���Rp��d��)i��&��_d��u)�r��MO
�d��:��<�2.���Lh�����-�<�6�T�������?��}���Q�|n'��GQ8��V=���ADQjĲ�R1 ���[���m�1�����KM_eʝ[��n�٢s���&���t����J��6���ߏ�f���E.^��$	f�I�xU������/Y/�(i�J�l���#�xG�B�/��dq,<MtKK`����$R�:Qq"�T���t���v���C��7��z�}P"Y����o
�Jh�����OM~�R_�U�UZ�Һ.^.3�rk'�l:�u�� �_��:�q�eo�)9�~�����yGW�ikJh��Z
�M�L�-/ʥX�.�[��ʢ���p�W#H��F=��9w���������Gs��b�\�����}�П[ۨ꼊|!�)�W�&�ѣ#'��h3�)�VU�W#�y҆�d�i�|p�w��|�&��}��N�r�
��,C���rQR&�`��Sq��y��2K�x��>m`�E�}�Ebt����I��K��w�r���\^)(%��y2i��;&d���sS���!Dۄ�|�[� ����ݖB-�P�=&@�N�"�}�����`�ܚ�y�7�L�a����.�������%�V��(k�I�:PU	*j��?���̷�a��ܫ]�=�~f��<YmlޡX�����(�.qD Tj�U��.��+e�^D�45�׷�sd9b��!ER�z�`L�љ蠩r3Q%��.��0:��
J	Y�A�F�G���l 5O1d��O�������nG�IW4K��f<���V�-�o ;o�~������p�"heERF��E��Z� �L�2F���/���b5�l*5y�U�����[Ǐ�����ӵB9�^[�]�uR��Ng�4|�M$�x;�ܦ��?��t��<B��5�c.r���8�܍ݥ�t����$Bϴ�ݣ4��l!\r
b@[a�1�K킦���	��z�!�:Y-%�Wu�ТU��$e��F3ξ8cm=��_ɶ�̪��|蓫�[q<����꽕�N���Z��T��Un�B�urL�̢�t3c�(�%Y���( ��ό�z�^	=�TM���D���"���s��hp��}����ۗ7S��3s�v�p���o��&z��:�G�����h0��(�A&������Ta"�V��]#�g�Np7�V�����g���C�Ƚ�*��4���H�Zϡ�D�0V(�v�����(���'sΪ�V�p¿�\����|�U����[�ԼBFe~L���A�1t��.�L���L������5�Vd[�~���_��S>FV �,�}�v7������c�:������b�e嫇XCT��$��$u����Ծ`���*��&��O����0���*�XX`�!�\�|dW����Ppۀ�˄�w�m�&):��-~Ǖ�g�͢#��z8��G�:f{"��I�0���q�s;���a�-���puL����F(��}-J.=���V���-e�,$�����f �W����E����/{VC>�ğ���[BԨuΛ;v�x���� l��?7�ӫ�ň�� ��<1��(�}���/�VK 5��"
硪'�J�Ӵ9o�Z7o1_$��#x݊��M��e;h��������>�W��s&�찙2��ech���Z�V|����2AF����Jh�����=K܃�24���o)����*6-`���/�v�W�%,؇�������/�i:_�!0轷����XG�6��3��w)ĤBS���XK
Q�6R�RJf�,3']���J�w�Yo�f�J��6�s9|��Y�Y2�v�o1	{P['�w��)�?˪n�%Ʈ�5�Q2��nP��N�%���=�
 ��h�~�������̸2'������$��K �3wͼ�64��Z�Tr���=�ŝ�CB�4�`�RüM�r�@��X�.7Y{��@,�yfw�VZ5V�S� �c~�l��> ;�y��L�(�)%S����RbiZ�� �uO��/�V��R����z9��ι�k��Ⱦ�X)�<�@K(M��řV�aɔ�����t�M���2�;�_I���x�p�ݎm$NY��[1�.75��q)��J	䲹\5� ��mag�J�R}4���k@y����O��ll�ԛ˰��w���4�8�}��@�L�_b��Y��)E���$�}���N�X9V]�$	/|ɑ���i�QL�}�Z��_Gx:�4Q�WRUb[��!r�'��[�#1>�$�h�hH5s'T&���{&V�# ��+��2r>�~�L�ݒ���m��OT�7�Xp���n��o��^\gD1u����K�'"/�:g��V���=|G>�X�@�g|��+s�ƕ�����Z��:�%[�9��v�"{J
W���=��s��8�bMۺ�w���x�(��B��*X}z�*�6�#��	��Da9���W�8���"0G\h��H�mrV�lgv�������GU&�ƌ?�+ޏ�[�e\�L"�UNDp;��x�pa;���fi�Z(:R��k�kI��bX�aD�0�H�w��^Xk�HR�,�m������ �����$;V	���"��]�z΍lm����W��,��ʴ`ܸ�?츚uF�嶇G.~�zb��T��A��En)�tH�W63��ۢ�]�H2�UM�%�]�Jw����|=%�[/�6�Y��tFq�59%��B����Ȧ�X̫I�[W<'���B���1`�xPV��H�s�N�����|}5�d��`��=Ϡ�V�������\ۆS��x��`ܢj�!ٺ���K���*G�IteliG/H�@��{܅�=r�<��oGZT#�VL'Y��v���E����p�=K�����N��R�.�D��m�ű�,���ԭ�����H�хqf�2���0:��.����VU2>�%�H��Gh�a[�&�k7�ή�ecy�:_V�2{)B����� ��	�ܼ���1	�N_��!%�&��x�7���4��B;)b�08oee�B�x�ӓ'E٢����Ɇ���KgݘK�	� ���~����K��H����|�;���(MIr�+�kd���"��2�uȩ����=8I_���X���W+��r�b��ڥ�h0��E�,��9!N{���Ri} V�&�mZ�~�p���A���
�H�0';��[2���ݱ΍��
�É�F��1�[8����`��bҭ��������}t��m��^(�/
�JM�L\�!�u������Y���2$ �#�b����a�)/�� �t}چ��_u4(�Nd�)|���;p}+������e�y�\;��{3�͹(��;X��3�j���2�=ݷ�!C�M�V�I=3ju��Kةhvp�b>���1< Vß�$<�JTuH�5�~\�
���j����i�kq���@�*�3��'���-�S}( �8"�v��>�O�;������h�#TL�N��h4�"K�b�����Pʒ�k��B�s�#�����e��^�Se���$#Z#)��N�ׇ�L� �iF)uMF���q�L��/ج所��e��wO�e3w��`��{'�D#j턒U�Q�yoϋ9%t����%A6������ya�`�M[�cWч�I�W����"���~	K�/�(�|)rx�6�3�W��#��gI�`"<�u� `V��*�C�S�5�ν�0��^��>�8H4G�N�PF�f�R�L\ �Sњ<)�AH�>����,% ���2��5��JkL��7�7إQ��}=k:�a$�,�ibQm�ZSge����)A�c<NP�1�k��z @jK��`؅�,�nq��xB�o�/:5W):�ڼ8���q@����vU�L�q+������,�s��K��Oq��7�ʬ�l�eٍ|���,�eG�A@���> �7���)���Z9{�DQ
y�Ң0bh��շ �OL����ꨩ��;��s[
���xC͏��Jat�vݞ���Z� ��t
	��F3<�b� ���)f���'�n��t�R�c{R� ��5��������[3p��.��'��=w�.H��e��9.s��Od�]�^$��~�K��H�@^%���"�IV��Q���B�J8c���A��`�⎱�hn��Qq�R
:�ֺ�	m���Ѹ� }È�A��_h�=�E1���� ����p�OuH��l�i 6�|pھ���Zh'"u��~���Q���T73�s���h?O�����۩��9��S������i�aj�A���k��7��%�5r� }���߃
x��b5�*sV�]S/�,����*U ����ֶH&�$;��G
�v��L6��:���!�R�AiV��t��z���?!�l��IeA���U<}d^��=��+��>�Yrl�\ۊ{
<�q��D��X��_�Ѓ�&]�6 �i�5��_E��4"����Fh'G���c��AX������;�N��0��(�R�"�Fq8�לAD:�OkH��ų�@5{�F�6C�,Sp���\�D��W����A$�4��ۙ��aX,L._p�'�s���6��T�u	.��@���?��I��V򿀯�d�o-���ŽP޷Nb�����n��6�=0VB�$O��A���lS��;[V�E@X�x�
(��.��k	�:�t�m�] ��f~;l�e�����%6�ڜ��k^�F&��H7��Ѡ�"��v�؈��Gz�I����F��Q_��zı��7cr��VX�k��@B2)F µ;�����oiN*N�휞R��-ˣ���dnʘr[Y���� '}��-4e�a���U����<ɀ�7ŐΛ���z�Su��Q�� {u�+�e�ӕ��rث������72� ��E�q"�u��.v�<f��]�?�>5�O[z��P�" �u�D��ev�=kH�|� �����'*���~���,�(O�ϔ>ku��&���b].�z9fM����mӐe�Yp��-Kw��h�b	R����;U@�b�Y�ɝ=�72���G�\!X-b���rҦ�5�� ʎ�6��> �� �����_��D.�X�&�A��1�]X��e����'b�'�N��H�}�[,8R�X�� ���������:�6��1Cڅ&\�ḗd�GC����*eO5��gF�[�_nEnC����v���RaEu�$�s������Q��IJ$�<O�b�
H��EG�RF[)cX���oB��}�<A&�h���V�ܟE���]D�V��]g����jt���;�'��	��άeߗ�BS��Oh�(d�%s���t<a�)��Q`C@�|��%�:�7�)LpY*<�,5V�W���7h���S�c����{�?�\me�����m9W;�cw�u�o��������) �:�i�B�=X�ڡHh�`|}g�#��О|�RA�JR!.���%Z!2�c�EZ��Lsh��9�MW� �T�mԘe�������GNv�6ޔ���f{OɘA��]���'?��_�H�Hl�2=:SX��~�K�9�P����{y`fќ��c̘N��P6W	�n�E������+h��Zs���%۾rb�:̓MW�r�0$����?%���$�݊��N���g
؇]A��^"�w�x��S����m�c7��G��M��o�'&#Q��%�5@�N�m�S�h5�]O�C()�/���]��r��Ʉ��/M�����o2�s��o2�����ί.�Ԕ}���Z���G����K�K�j��_~_ޣ��BQ�}fhNVL�ߴ�-6��N�{�W�4�-�N+5�|4_F���:����Ŵz>H��TI*�<%{9��1�T�
�B,",����AF���� ��٬w�"�ը7��?Vd�,�'40�<�³���Ё���UV�U�%�����D��HE��$��g��1� r�t](���}� �0�2��ʱ�%���K���N�wfu �RK�E�Pv�����D}R}`�m�q��<���  {����`�]��f8;���W�T�BK., {��U��Z���(�[�苫�c,���´��w�owL�9^qʓ�ز�c8a0�^M1ϳf�>˖��ɳ�y��}]�O�G��NeZ�![�]J�M�6�����������[��em��͗Y���a�"��!��;0�֣�*�C���L�����s������?iYf��=�`�s�|��k���~��pD�Z5(e��s�Y���o���E���;��L���յ�� (ҵ��NY��m���ַ�)�}�zpW�x���[P��ڕ�acv�H 2��!ӧ��̨�k�b�o,/�����_7�{�����c��;EP�"
0��i�.���������7W���2=
�}��$3}R���L��5o�-�H��t�:�kb�sz�zsV7O�(�\��N&��L�g�)Y����/˪�8N�˹"Q_	�3)���/m�	�a���_6/L�I�p	�N'�����ɵJ��o�=h�{�����|V�r~�A�ϫq_��ӷqK��b@t�1r$9ٹ��D��6U��U:\(�N�u��O|��L[��W���ef���!r�B�z���gW��Y�i��p��;B����ٿ��,�u��fs��Qv9�P�E�';'c!"'��wxd�[JO��YՊ$������/��ò��nb�%v�
'�1�;O.ugz{W����}��h�V�Lu����'Z��r�:�B�ؔ,�-K����T�Ǯlױ���'��?�WĒ}M�^��%$�-�+�R���,����b�_Z�Z��kɬ��Koӿyp��:a�a�GC��soE�ep7�`+��Pۣ��=p_o,�������Aڼ�k&Qc'�5L2�6�d�^U�[w���y�@3Jg)N���R�y �i�R]Q;����^\�%�I��A��W��Va�x8��w�'RO�Hh4����Y�a��츝�9�ހ ��	>_J矐��q�����ID5��{+���m����HU�6W��7K"S�GAZk%�i�b�ay����g���(3T�bE?�"b�v�)�P<X��;���d{r��R����H}�A����.�2c��D��(�G��;F����.p�爛��g���|��8y{̖"�t�9�����}0P?������.(�kR�D\V��+/�������wE��NG�Ѷ��/������AV�;q%Q�X�	�gb�g�ls<
�t�G�a�w�T
	
_�������7��e-��cX�6���F1fe�#�lݙkMٞF��(`K�lZx��=�'�+6%��ўZ"i�2pWQ��2���n�w��M2n��Vjyu/^��_3��]���]��	�N����E�el�3j���{�,e&�Z�a� #�W�S-��hG���+O	5� &3)[��T����LM�a�uK*%1�a��:�z�ʈ�s���x�\��9_ ��r�������&Lf�ȉ̴F�-ҡgs�����i��Ԃ�S����k�K��BM�C]/M�@;$��[ �3SY�C9��&�2gL��R��T�`*�SX�zm�� �W�u�ڿ%�q�Fzț��ݝE�]��k��n�P�b��8�t3���.rK]�.4*���щ��ܿ��`�]���v��O���~�s&��鳞.�[P'�tf F?�^C#��U��]����1����PR�qD`�|�I(��߽s��<���Q`���<}�3T�_��_�M���-0Ѡ����!PD&���R�u��3�0�-PDy����<u;���ϔ��e��S|�,Ԍ+�Xi�5�%��&�����IS�>J��:D�F��ob�������N;é%l�t���|��]@gߚ��3�H��~/��{���ZOv=���Fd@���DG�J�n��]��/Q���Y��=FS�[���ET;�<�� @Z������Q��c��4oh{Ƒ.��ׅt2��3R���\6�}��*��:t����ӂ"K�0�*�O>u� V�\���Sad���� ��xߍC+���Sl��1?��]�46�@�B Q�Nq� 9�^�*qO��;ޔd0tDN}Y�u �ԡ�6�|B�"�8 Yq�}W<���zb�)���g�Rx��E�K�D��Ԡ� _���'�U>�:w'eFe�&όwM���^�i�7��Z�۬˧�_�}�N?O�A[^^�\�c�6�p����B�b�*�3����|0t.kμ،������h�Q�jE9� c5���`��i�%�Y)�*��6e3Z�؞e�H*ˌW�K����]1�X�p�ʎ�� B�B"��NWL��ު
'��"%|�
5����}r~�M��Nk�$ߴf7T��G�ǳ۸�u-�(v:��b%�F۷d��8P�U��5�<��۸pޒp�����;�ʤ�}!vGҢ�]��u^ �}m)zQem=�G���2V�n��67bsRAPU��):f	��}S���G>�nG�g�5��cū1T/$�N�$!J�Բjʚ�n��ȝ���Ѣ�/c�Ӌy�ܟ
k�V��� �7vtw�W�<�˗���E�C�%r%��� �$Z1Ѭ�W�M��v���U���{��A����8�_n_ ��qzS��=i\�������'{x1_hȜs�|��v>��I���e=�yRh�OU|��p1W@+���fv#A}o�N�t���ӹ�k|b�'�>7�������>���y�8H
}̻�K�����de7�x�^��������$��^��$c��#�l-��-���s�g�}U���D�:��~I�ֳ+O�b|r�SO8��F}�v�3�<�y�v��ݯ(g6�߷'�4�^,����j��?�󜗔O�Y/�J���!��#�S�b��{�������Ⱥ�A��ǝE�V��R�O�u��|���B�y���9Q5LW����v����hƙ}�1�9h���N#�	��,��W1eTy3,���?)!͓�e�)p떣,��:5l�'�ৠl'��g�G<�.�i������J�J�! JcTQ�E���#"��V6�_��Ij��z��\���tv�	��n��z�����5�r="墲�-W�C�+s�.YH�/�Ϗ��*�WC%$�����
�PJ�hB��d��	/u�x�~n�,HxM5/cQ����_�XO�
�D�+�C�ݫ��=xF�-�����7J��$X�✱RCw��w� �AE�HVwZ��};P���m�W�J?�"~�|���w�wTX�F�	ڵ]�t�	�������uQ,���J����*�vu���|RV��>&��TE�hL|IM�JtM�?x�Z�b���b�5q�^�����xm������'r���&g��2�`U$q��˶�"D$&kTrt���`���T������?��r^�`6��a�$t~}�6�w�6�i�����V�Ͳ�$I(B���R��;���ï��Њ9��<ҭ���|���s�+�D{���h�4�J��30$���]���m$?��a���8@�^x^Ʋa��Τ�c�)q_l��c�I��B�To����h���l~mj���?a@�v�*�w�����^�_�u�G���@o�k�͖�oo�1\����,Ţlw�}�{��0���Lcԫ�GN�,�l��[I�A���#�vB�hxN<r��=�������א06�i���.�5J�C� ���l~�w���W��:1�B�>��:��a�D)uD@7tU=�:��b�c����I\~XU��5�&@�<�[����w���ֲ�_(�cĊ��V�f�0c��]n.�?��J�� v�ꋾ�oFj�2�%!�������f4Q�W�/�ehC{``'Ь�z�~�nhY�[!n�;n���YAH���a��JX�k��Fe�۱IN&�x�PP��S�-�7�vҳ^6p�x�w���h�t�+��S� ��I�3I��HO�9��v�\��NU���MPYs�D��x��|�y��*f�y|���Ơc�qu���c#�w���(7$����A�}G!����FO�P@�)7(�[v�{e|�NYL܆�h��9�_���!:�{�.�*�S}=V�tu�a���,��J���U[f�yЊL<����^s�:�e���_]K�ն��GŘ�*�vr����n.|1��;�Ӌo�&ɋ�O�K�c�Ѕ+�J'���D������ϧ�h������x�J���B�p�	��s�sP�`9�j⚢i,�ߡPs�&ޤ?�(���':^ª���w��tA��X�`ol�C惡�as���U��J�4��θ��lɟ9$��Cf\�]�O�:1++���WϹ���{Ya]ҁ���P�]��~.�2�xƥ��[�G�oMdX�������2'-j�g��4-��Vu	.��a��b�Q�a�9����p���)�����L�٢-{=&��4�(&�?q�N��n �J�f�P����u��A.l��hd���/�Y��2a�6�Х9�@&�;
�����Dƿ��ֶ!��Uid~�� ���ʌx�F1ź���	8]�[��M�4��Ga�q�?���s���y���� �ο��C����e��
�2��Jw��F�ښ�9zt�jچ�/��^ ���YE�UU��+�������h2{���;t+���-5?���Y�8�fS�r����-տeL�^���ه_�n&A΄`� ����!$ ���{ۯ9�\��6��O�v���&�.�|�d�h_Ԩ�T2Į>�)4�������? �]�}��@����F�H�r��ZsR��{��ࢃ�t[0��ַl�`(E�8H�t��\P�OB��9����h��698ž&��,���=���Z��RK7��]N �g`�k9�ň:��)�jrmQw�Q֜�����Q:���/X}4��ψI��g����ۦ��.db nx�)�R:�?hJ�m���t���$�����?��N�)����P�c|t"�{M�o0��ɝ�4�a��Eקлa�ѝ�|gǎ���Z��T2˟�q��?�v�a����M��jC Qq��}����J�'3�F�:�a%���1M�LR��4N�|�Cc֧�.ԙ;AWJ"��t_���=d���g}P���ZB�[F+�BSA�Ct3_�p-�u�m*7���+��6���d�SU�:Ӈټ!�H���_T�O���d��yDmcOL���L���ua�^ig�k��PL�d^GTl#L����Ҹv��4Q]5M��֣e7.��D�8Tl8n��7�=<9�8/�	���oO���b�*��Epʞ��V�M�'f�� w���#q�Ck�a���#Lݾ�Q�x��Y㎀`I� ��w�N̑�z܉XP	���,���H�7c��CcW<�?c��,2� 2��v�!{�����![&�Y|�ߣ�R1n��x����,��j���؅��겼q�B���5�p��q}�x��,"������޼p��>!_���"���^��9���-�Yk��Kn�i�u���O��E�GoN��EY��Q,܆��D;�7��g��~����.�""��U���mH�-�S�1<){�������c��S�O/FB��(��Pc�lCE��6�G@�w�S�-��p�t�����f����mX�[�k[#�tԉ�����4�)��*�~�}<y-��n�b�*����A���6�98w~7�^x2��dy��?
��O�$�%}2��;YX��tD�h�����d�2���b��ܡe�v+uafCOK*�[�$���_�������"EfӖ��e�mqdy�����)ϼ�2N��1C�j��6�>y$�Ji>���FYO�njXS�q�C�χ�ܸqq+�G\ 9G\�/�M�L�<��H-�6��ˡ����RO��P�n<�'������v��8����-%���D`��^m�)v��ŇTC��O!�K3�!��f�S������enP��n����$����0C=W
�<��dF8�qU^�ߩ���	'L��������[O�$�^7�� ������J��_����FE���.��%�sM�AK�}{�w��Ǻ-��S�2�|C8$RM=qtT--HK�I���a��r�(��]�d�D),,���+�����1Vk<Fry�#�O�"�{6Xi��������=�;��t��Di���`�XS��=�^����lw�Z���6��}���H���)��f3U:��c����wɘ6W~���'d1ބ�����!�m|���J�yJ'kW��9�jM�ss�)
�,����ݷBE�8Do�s��e��V˕%^Y����9�a���ޯH�څt�=<�#O�=�. CFxy��^{&r��T���'F��a$}s;����]�ȻEe��5b�o��u�?���|o�k��m�K��s�&�?�k�����G��ٞ&��FY;{m�;6���2�Vtq�����&��t0Zy}s��E��Ά����ͪ��+/���4h7��U�~��96E&����Z�u�?Խ����-z��i�Ӷ����P�1~3��zz�;���ϓ9i��� �f*���K5����qJ�䩻X�`� k�i�+ ���Z�l���?'}�3g���G)Ø��X����Z!������	I,�.@�P	�؀��9�AJQ���z������[����e�ڋ	1���fxQ�͎tS�K(�����	��R ?�z�7�|�#����[͹�'���7����Lr&j  (�)����f�y��O��沽����W|���2)-B��"�5�WV�D_ؕPTs�iX�?��pn��+$er��&C_���N��Y���׿l�Ss^����a����o�m����+9hL�/��^����t�ʓ	V�܃!%x�����f�f�����aͺ!�B�RN{�?��9��Ӈ?A|{P*�w@����	8ĉ\���z)d���Km����M�-�ӏ������r�d����fhO����D��@%�+ӏ�«K�����{*QI
�H�1/:���?���]m/�x�O?�+�����e�]x�W� ��}�0σJ��r����"y����]�@��Z�D@�&/�ŠB��BG:�^x\��;?ܙ��\�A���Wvg��E1��◓��K��N�M	�*-��S�0�E3�:�J��rx5���>1�o����VL�Ӡ�����vbp��?�|����ex����N������$3��d�y�y455	Ʊ��V�Q���atxգGI__ ӫWOHYh4Ϳ��\\�\eQ�d�؛c.y:��f!�=�G�hl Y@Оgk��7�t4�b�i$ƣ	]�gvb����t�uG����������X1J8�a��A�3�T���DE�����]�?��q�%�9��CI�R����y_=/P�ѱ��RS���m�����35������-)�1˴T����=]ʄ.m�v�Nu�R�����Ϊ)O�)�>���/>�@��M�����\M-%9��7�`��"��}M�U�TtD�̿�gd�6'���j�����@�\~%�5��'7
�u^��>@PH���7�j�5s��O\攈r=ϕ#�3��Ǧ�{
	%�Pܹ 8����uR:����Z*��e��h�Ώ�N�M~�.�ь��T����A�F��n8�0���[�	g�%HXǮ�*�r�"��wv-dȺ.����$��gBm;�9��Ov���S�QA��:eT��\:	�,�:�N*��a!�J����9Ъ���C!�-<���D�/�i�D|�^�&ZEh�c���b���tnX '�ؔc��h�w��;�J4���
��	�?��T�~L�K�:bN�s��mТ�^,0��	cy��Z��YH�͉�L����s��T��a�}����bH�qrq���cue�G���o$�X/)��Ut�r���V��`/#��r��b�{��y?'��7b�X��G�bB}�s�Uph��觶��D^Z�M3ʨ0��bq���WVZ?Ҩ����ޤ�1��'�j�O�����d��Z�o..�
�:�6j�q��v�0�hJ����֬F>���_n�q�D)�(^ɀ&�Jr�'�^���� 0O��nS5��딫Op�Fpf�ǚ^1�<B��B������v��9�#7q� �����Hvlܣ�ŷR ���GJY�����y���ܾ� ��R�P��O<ӷ{��,���q��������m q^��)k���W��HK��@���H].���;�s�tǟ���$Y�k�J�z�&�?�V�ޭ�M��h�gA[
���Bn3�&!��{���I=z͉��O*���㹔������e��W3LB�Ba�ƣt۸�I�X>�*ի�M��I�`"���1��s�τm���<(���ZM
�K�4���&��;*�mݱh��5��1�)&,�//'�<�Z��X����dG����1DًVT|�k��l���3���i@����U�q=b��}z��5/��-kT7���4��3�`_���{��AC�,1x*�@d���@��T��3Ykr4�:���]��i��Zm�N^���r��B�R�SY��)ϟ$6ׂ�	�I�f��)�\+C�Mְ�4�9�w-�f��h�Lf���SA�q�%w ���X/��nX�H��偖ˋ
�g��o!�2�&���T=n)��������vT>��p�7%GS����/�SJ�������^ir(m�@I��h	< �R}�C)���F;=2�r��V�3�hѫ]�ŭ�w��]�{���/ŧC��-�u9�	��J���#C���Xcr��{C0���6�$���.�P���7��W"{g<��?r.��9IN�{�7!���	�nA��� ����t���E�\�fQ^�mG���`6�JqN������Y)v�z�2�>�s��N�:O`aQ��s����"�j�����WkɎ�1�iKf��ֽ���o�)/����'�(tҨw�8��s��Nj)���`;M��0���%�����:]�I8��cl`�:ɺ-����>��9�P�Xcd�:�sű�[r�y�z
9��E�����L|�#�R	)�����|�FfT��[,]Бj7ޜk����yv\Z"ְ��3���Xj��+�h1��4V_���&�d
{ɑ�!�����9�;�[.e.:�̗�y�.�4NT�f��#�д�G:� S�y�}����3]�3l���&�ͻ~�F'w�WN���W4X=k�p�77�62�M��L�B~�फ��������i��Q�Z�h|��<=蒋�NE�S�ƆSj2Ec���0���1��X��𩪟Hi�yFl��M*}���I�����jZE𫷜q�h�,�֞�1�H�!�+���&�/��m����d	-c�1}'�f: �s��,\��鸷��pD�^}Cf�_@��^�����<��'S��_E+���E��c�u��~��I�]���#U��+-�F0-�i�ȣ�E8���ވ �q�ä�:�%�IsR_y�Y�����^���il� �>_�j��K3�����{���H�_�t��S��A-��Ʋ0����U`�ޘp�A���E�#��Tu����'�<�s�ߒ�'Fc��c�͕;��X��3�ش�l�.3cmZ�A���R���a�(HL�"D�R~��5�핼�!���L��1zi�r=
� %Z�""$t[��4���3��
������	����9i'J5�l�1�p�2�|!"5�ЄP��)��N(�E_��3&�\2T��B�	���_'����;H�K�q��M:AL}�2t�c7�6���)�B�|�7qG%>���Z$~���`&���?]��
����P;&�f���=����/$: �J
�E��m:�Fԫ�� !CE$7J�l�|�}J��B�m����"����=S���r��Y�+i�~g`�O�ㄚ��	[�����B/;{�Ag6�;{�?�;�J\J���2sG��y�<�0��v���=�8�W�-?��V2R�����__V����͡�^�S�������es���7�����I�̮"?�[��������ڜ�^�q�娧PTjzj�o~O�i:�2�H7�؁�N��]OԬ��;��6��-���Xr];�2x�t|���Q5_�K�$B��� M���y��3�p7��q����y6qx�*.�
8gU�4��:�@h��Fb��'S��vI�|��PV��p���
��.���ޏ��w�0�)�ː���zU9S.O�%�'x�q�*��!�^��ڗ�hˀ�m?��w��?u���^�|o��S�+˥do}��{մ�>x�J�E��-ٗ��14�ϻ�Y��*ɔ���V�A�*%mn�I@Y�H�8a�f'�d��f�)�5�
���ɺ�	A��s7n_��I4��[�$[��������t��$����y��.i L����O�~P�l]��ٌ��=�)�o����#Qc-�'c�6�`~,��g[�e��2(�Z�+�V��FZSevڳ[�,[�Z���<���3��SW�Aq��n���Kk�µ3�
ZGr �da��vA�5t5��<�q��c�s��2|ÍLA�B1�^�i���!-�z�k������[�}�t�J$�Y�a�a��ʢ��5����渒+��#
8�9��叩´-�n �Q-YB:RzKu��cjP'�瘈�f�G6;"2#���]�`�/����=��WZ�/�ٯ4�Ҭ�Us��3)�������&�A�l��>��N�i��:����N�)���	���ǖ�1h�ھ4F'N�RR�D%Z�]��ȴ���ɏ:���ޘAr���d�T';@���-�9�뫊�z-�B��"yN���V����Y������(*V�f��S��Uz���3L�S��<G$�a'!ߏ$��IW����e��K@�Dh7���0�I��~��g�wȝ�\K�s5P��-��H�a��l12����(�ЇyC'�*ʑm�*;�����rIV=�� ����>��F)_�S,��X�-СJCo$#�a��u~A��Z�~�Z�bTЍ���8�*�����5vf�� ���e���f��%ģ�-�RuH�Gn�����Z�6Ӓ(_;���g�k�._������&�(4���Y�ύֈ�3������7�=��ҝ�Ə"S�+�+1�FQ�X8��Y�ѵ�	R��c25
{����
�Y6Nl��up,A�h�}�w�j�ub͎;�?��Ĕ�S6>(cP��4��}�hIK��Y.��^�AKd��*�ᷗ���,�"uz?��<ye�@p�7�oR�@D�^ M8CL�%���׃��7.WK���l� XC�����B�ʅa	�^e�����
`;n�g2���7&����� !����?a�;aۅn��e8}݋-z~�>'pr��znaua��h�h��D<�u���Z��3kUdX��44[��OA`Ur�s�h�T٘]i�-5p����\ϵ�Dњ�-:���ui�XL&��J�_�	��W�{K��. �D����ps�P8x]�)2|[�G)��$ҥ�;.�m{����'\�έ�Y�Wk�'�i?�!���	+��:%�����|e0"�Jk.�&'�t���������+���v!W��f���V��!��xj.�:�Pk�ܮ�QFS綈����rU�a�9]��^BYP:U ���! P#J<����W�<;�2�.A+��5��%Tek/�~@��nf����䪋.��j����J���L����5�Q���Ƙ�E)IOzv,F�&����/�yI/�v�B�
%������Phc��gĥy�:��H�fNdq�W4,�?�Ԗ��y�wC�[�״�2�!�5{Lk���Ee��	�^�*�V(PD��W8����q����>#wyyx��ד��{L�l����jZe�k���0'�l	�{`ǆ츍v�5�ql
ZE�B��{�r �Z=�����A��<I���HG7�V�tS���}����9jU���	�t	qF����&�����yb���ߋ��T`�U��g~��畋����T����p4�;�z��b�X>��EC� <���$����;Y+�H����5��,�7f`�����:rU�6�䀴X���	)����ԁ��r�h ���yRC)�\&5���:f�;�M��D�KH�Ȥ$��-�ˠ��Z��j<��z�d̈n,��gU	V��Ԁ�p���ǲ��06����/Gt�
� gj��7 �z��)�k�A�L�؎쑣d�ǟ�9�`�1A��-R�1}zʲe���M��ӥWǃW!��΅���Qh�^̥xh�Ӆiuhv�<�c��]�g� ��F/n�����[Ͷk���)�7n�wSZ��p����H��]�~��;B���ašo���9I
�}Ym]�LP*��(q�@�S���(�Ɔ�X�K�Sn�/+�?(n��n�Ɠ@E<�dgZ{���G������CN�hQ��t˞{��Z���)IʉG(c�3�g|�G�@�bf�ޖ��Nq���&q,5DsԆ�(<u���e�uorCQ�a7un?`KL�W��n�.)0��|��|b�N�]���,��<�18ɮ�]���E6�n��3�`!S�A���(�ֹ����];�����|�҆I����9\���ة}-����#����8�h�a�C^��c����H����or8�A����h�K�ә�h�6��\�q�$T|IÈ�% ����{V�C�*sӕ�&~")�e��&4�!�*�Z��؅t��}ϋ�A^�G�IQ�!I�$:�7?1��6��QFt�.��8������0��15�+Lip{�$�m �H���u����tńJ�{\�T.y�L:����./^a��Rh{WN�h�V���)��/�5�9�7��j���@�1��ڷ�6���(_���k���)������3:��9�qw�Ǝ�j�����Ч^JP�Z���<v[4���(UF�{����vo���Ӕ��=M�:=o��y)h�s���°)��a���G�J&b�S�F�!l"��	�73r�1:�P�z6���Q��iW*��y��D�,��o�:u��p|�'y��9f�[Ӿ�� Kx���;�;BuaC��`M_��xu�s�y�m��M?-�����CS��̆�1f؅�+�8 ����%ݴ,�]���Ϝ̇���L��{d�{N��f��Y����XN�S�����b�����S�H��׈C�UCO
�\�y����[�~#��I��U	��K��J��l��I��݂�~���˝��)#C������C��+���&��y����	 ��W.���V��x���$,�Z<.��}/��`;������kƜ(��VE� �`\(Z'I	� �Z˃��p�e9�P��Y�׺t�1Y$�`�v��+$��4B|����Ն�1G�4����Qs�t��\�����#�@�����f��njʱ��`ZX=������j%�`�Z��>�53E�Nn�ŻkgmT�v�`-���]�*�зd(�n.����ӍXP,��3�wt�>�vAc�7���cD��q�T�KG��1��p�^��?֒0c��DZ:�h���r7	_Ғ��#�2��H�^�a��[U�I9��m{�R�M\�bO9 /b5�UJbG�'k򣈴]�@wD�GD�nNOh�I6I�T_��~W���f���V�0~4P=O�YTV�������
�f2J2��|��~�R7k0NjDx���S���{��N�5聧.hLK�{��Zq�U�,���k��{΅��4޻���uj�=A	��La�״{	�}K�
t|�L����J@f�1�:���h�����e��0��)a�>֛�f�	���Ϗݛ���^;���4��B?����ןS����8��A�ɾ���9f�y7MJ5G��@W��zi\��W��;L�xE���o21�ӑwe_�O"nn�־�M%K�~�my�~�hݒ�e�k]�p/}�@��`O2B�b��煇k����N1���Ơ�]��ĊJ���b+��4�*Gs��"�}#�����Yw,\���ۥ]�c�(|���N-�'-پ`���u��Փ�(]��c����+��o����p�W�d& 'Q�cL\�~~Ȭ8OL�՜�ja�,V`�c&1�F�lU�q��\
��9�R(b�N��i-��m�̹���T�K�.N|wh���,���+#3>r����ߧ�HNT�Q=���| R�Ys,8���p�-�y�&Q�mST�ت�9�V�Ur��砣��I+4�*ap����H�K���W�����������>gz��S�X�q�:|4���D��1�Z��ƖFy�pj�]��e��+�|r�����,��W�=��7�ᅠ��<�2��I�i)E� ������o/�g�V���S�i��������>��{��$�%���)sp�XTk;)�l�!J�.�+gm���"�5��ߺ��Q�:V� ����п����p�Q{�Z�cར;��O��8^�8�����D5 �H�N��Lӄ�d|��3x��:��yh� +� �9�L����
�(���{�:f�T�����7�?���Q���Q(9�NH�#\ �₰�$��7-����H��	@�T���ԛ?�6(��PD��(N�&�1����_= W�9���V��^O��E��ksU��.�& ��]���$�AZL� �s��'�|�ȇ���u>��٣�E�EA���q�ve�X�H�@,0��k�y�*<-��"Ȋ�S�9^Gu��g$��n��cU�Cr�p>O�fW�He����; q�PDV���8��|w	餳�C=�(\��j#v��Wj��+�g��|>�	<�$M,�o�<��ѿ��i��Չ-ʹ\z�f�xu�[�:�)�d�`1�r��Ǟ�Q�nZ�+�Wi�d�3̼+kn���)���$>p��m��t�귩��J�����/��'�)��̚�;Z1�NT�_ϹhC�dc�_�f�����@n��	�-@}��$�c���@���I�[9���䫱�ʭ�M��8�N(m��&����BG�=�(=D^q6�v���+��ʦ����A�<]������֎�{ƭ7nl�7n�a5�V��O��{f�~׀��{E�O��bX�o�sn�i�m���ի�6�C���_�'D�
7�l���LN�z>��.j�et@Ü#����'T0]��KW���RӠL�}����φ��B�ڙ����7��9��7�ȴ	���~u��rs!"s�<&�ehh�O���z�0B����@�v�=���dk"O��B���y��<T����x����[�Y�훻%���愹][��e*�6n]���0V0ń$E�dk���H�h��gyR
���y���kKLL����J*���.�n�Z�	�W�\A�z����KX@#�s(<;��4���F�9�A1-�d��d�a���o)��*��&,Fy)��:ʊ��=�hx�����w&K�a�*�X�o��%�(�3$���W�O�7N���x慼��>��#L|�jh<:lV�[DX��߸K�C��p�E�j�U{�3d߰r��=�Qغ$�g��2-z$��6�Y��_)�#�ix���Jwnƕ�bb������<���h�`o�Œ��� �5�^�M���X��N�es�[H�MDE%�5���U�cV�Em�r��R��=ӂ����?��r�����j�-w��I�Z��|zb�*j����~������6�5\��˷&�Z�����T��є�K���w����������q��G�ē�!,pW�8O�q��(Z.�r�cH�'Q��iҟj���	ve�,<u����yiw��plz��؅�u�n���~�e��ظ����%�"j84ۦOu�1��z��W	�,���`^�����ޛ�%��(_� l�AN-�����"�gu%� �
��J=�'2�o�ju�S� �|��,`]A�1�0=U�)L%�uۙ�%�B��z*5�D._���z[���"�'�������9N��M8�1��á2�r�{�*EE���țLj�=yx?x!���S>$�/V�*�n��5�w�W#����ݓ�‡��Y��[ٍ�'��!E}������ޱ�PX!�\�u9V�/��x!_�V�kg��ny[-��%�r�Yo���e��b��0��/`N�����ե: ��sӝ*iT��F�tC��V�����L�@����L2c�нEr��Ǧ^.la��%�&U��1��,"vxW�w��"��|���L�4��p�ޕM�B�5@���q2f)V8t��DQ��`��9�����)	MA�A2tܨ����Ɂy!GI��X��3�4����G_Iׂφ@%`\��[$�r�z/�O==C��7��!evlM @؋0Bs�� [uQp�h�f��o�S�goJ#.@py�r�v�;O�� �ym!"U� c.8�%1�,r��c�4mŞ������f���QH�	����B�F>�	)Cf�}ҽ��#���m��MD�_�P��>�����. ��:"3��8ނ��&Y�0��N���c���0���
�_�o	�� �ǉ	�����A
D��9��}��
��e�j�[~_�@�h���~���uﵨ>ΰu�#u��Z��O���y���,�z�C�@�Sut�-N������p�b{ٗ��7߾$fTq�)�3����e�䵯������v=�&�B��]�Ӹ�uT ����n9l���K�4b���8e,��tYO�R7؞sR�(� �et���7�[���0t�ܺ�K����RG��I��R��p�w��á�xE�b��x�>)�������^�I�
�mq�o��|��X`�+�s���R�~7�|[u�����$;�Z<�ＳP�R{&p���Z(�c�n���t�p�*�(Z��1��pJ�J4r�A�T�3n[�a�����rb\�.��mU6ML�e#��j2m��5�+ �H��+�s#�/��iLB�9�9�h����vZEzx��q������˭O4\O�61�	�:m���wp~��n�	-�JA��T��-�$�$YÁ��f N�R���e��B���(��ǌ݋"b�@7��Y�ׅ�h�j�7,�����"�s�()'D����b���ETe;�TR�����x �I���s5���R�1��)�S(hf#�L�Q,N�i5���v5Ld�R@���4p���%Bp$
��au�5aE�6�jS`ȡZ</kBC��Cܔэ��iI��ό���X�ޗFNk��@����J��'��<aJsi�7u.���LI�$����B9��V|�b�d�l�ʑ�}:�� �`2�S	/`��/�G��T����/cY/��[+�}�(ˡZn����B.��Q���$3�%{a�,B."C=(�C;�����ܛT(���\r�4T� ��m��!.���V�wՆ1ֶ�)$�L?
����ǹO�]w0���Y༊�� J�8Fᨋ�H�
�u�v��+�_o$��qV�q�������[��N� ��gٔ!�F�#v���vǆ��:+:��(ȿ���C�y�Wi/�x�p�����u]�"�fd��wQ(��~$��XA�f�Ž[-V$>���
��<���>���ޖ~l�e�uR���� �ys�l&��Y,V�������"���.v���'{��f�!�W.�M�Z�8	�ݚ�B~���A��!�5���>�i����ych��H��T/��s�H�������,��g��&�S	�@����f�g���;O��<����Wc�*��#;C�"I�����>��B�������C�+0�������$ĜKNȷ*�#1h�6��LP��_`���N�`#}D�%��GL썾�E�P�O�$%�������XDZ��|�]^z��AD��5ӽfw4>��߉�#��n\q$��fd�w�cL��&(A$�v�$�Gwx���݁U����V�L��]�u�8/� 	��}P6g����2�W�,6f�ݔuh���zf�,LY�{�b΢P��?�\�λ�% i4�_Xi�]~KZ���g-�T��p�������v��g�"0X����"��8N; �ǲ�Nr�)���jlOsr�Œ��g�޻6���"Le���$I;�=� ��1,-�'���<�`�7�C�=��l�C}ܐ�9����:|�d
����O 6��ʂ�����^�1�K!��":�޿Lf���_)�m`�9@�8��������SCNN�Q����N����RT�賮��f��O��;]�_����ITܥv��U�����\�`�6M����.���ƿ S��K,�+j婋�?3�������m���������ɗ6��$'][���{I����1Zy�m���ZmBd���S)D�����O�v��*�`�q�<�-�0���w��(F �bfF�r:��{m�b�hUf	�O�˽����/�H`HH�5�����`m�K)�����#��c����lT'���d��3��U�i�K ,�#���Z�@����z9��jMF2@��P�y}1�l(��Z\x0�7R�o(��V��
��Va�ݹ�&A��*?2��v>a�/ũw��Za�t&%��2hb;�V�VT�B"��� �!N�!��b�픔��9��?��Q����ٳ�J�;�;��Ә�c}o��f�)ɕ�����6����):�xiO ׽��O� ?OUO��Βuh�o��#��a��v:�
��[G	���*L7:{���/i];a��8�JzZ$w,����ܞ�V0^~��z�j��>�ī��}�7�폶��ȃgD,��;[ԝ.e�?h�v�������]d�t�Q�_���BK��$���B%K�FB��s�m}�B�A��g7>�gʟJ�ΥR����k��F[���&���ك���$jJ�U��k��͊�Kuҽ�_0Q�ע�d�hԓ�j�%�s����gbG��ƃ+�3wcx��3l+݄����?� t���C���U��Amǀ��.@9�e8��g�$�����NJ�/5��EɉH��VO���X�$�t�� p�0�7�_HD�����:�^���1�=�e��w�e������(D�o��T����Gb�?H�*�U�t��g��N���I �=���e]�,��0U����n��)t��U�j�F����\�<s��p����Ʒ3<P�X/Y)]���R���W%�'m�>���'��guUE���ይH���]������e�9苺õ*��Bԣ��b�_o�[�7��c�8+���$�(��@j��gf�lP�����6��N�N$�F�X���C$-���'� �^7�o�W�r�mml��|!�a�lX2@�η>ѱ`�:�\�a�R~�]z�ũ16��#B���p��:}6�W�ҟ���hW\r}�|�@�"��M��:V�ߥ�ge�ty�j�sb'��
j�������%c���)�C6�u�4�4�X����ysq�u	q8�;Rk�I?��p���9	,Bj��X�Q�%� �v����#p�3��>v���� �I6n�>V���$|]�����^��>M����@�;�����	~�\r�E��j��~�T�?D�w
Fx1_���M;��������O����h�{�M�1����B{+�0ri��6�y�!���~�kH[�ѡ^J�2��	BErPmG,�7����-	�-�wL_�M�`[��l˨��>-�I�N']�PW.ǝ%�j��޽��)so�/�oCxt��i{���Y"w����p8cF�D��_=�X�D,)�K���kIШ�<z���W!~�+���n�P�b�u�؄�r&q�V��%�$U�E���3� !i�G�o���>D�2������0��%��ܐ������X˱�O���6�����,��	k,Eg��F\�ƀ�͜zB�<�|@�ڻ��F�������4����֏Ǿ�!�����䖗�;{]��YD���b!��!����N0����Dv��bw��j�S��<��*Ҡ�I0G�?�M�duO� ��\�e�����?��Wz҅p�Y�Eiw��^0��1��z@���r�v�a����Ҟb@����@����Oqm����W6�$4:�����8��\!����A�~_��]�S�T��)# ����M��1ɶ؜���Xa����o{�����m�:�F�Y� u���|_����?R:^��]�+�k#�� ��hO�!��c=�0�t1%)���ǐ�Pm$vБ"���t��ڇ�Bl]dZ��Rq�&<���Rb&���|ՙK��@kNBRa}8n�ę�Zu��x��R<ǒ[��_��:�m��Q\��F�`�?�{r�@������u���3�.��c��O+d���;�
-�u�;c��%XM�Y�uY�o�<�F�rI����!����ht`.���@�m׈08���y}�D\�)ߜ8?P&��<��2�T�s�U�B�%�Bײ����Uam#��w��f=�M��F�)cƆw��¢�4���O�L������M�!�-�h����s�"4!^�T����w�M{<<�[U����4�@��*��6�;q�J��]�
8v%�=����j�������_���vw�����};S<8�Z-�	*�Ɩ_��g�b�9�6��_�~�|ϳ�Cn~G oh1rI�w]FZ�ؖ�������܀�C�jkvɭV��(�=�&J���qnY�Z���s�����BUw�t�n�|�y獮���<�6Al����B~V���6��?E\�e `C�ȳ��z7 4���V��h��1���;�39E#3VV���s��_�]�P��"�.v�E߹�vC������_x9G~����'VF�M�}����n��
s����d�ZN,�R���#�u��nZ5���bJx'R�2q.b5	XOE��E�Z�>��F�d��춄h�S�;�J���ǎ�F���Lh��F���U��>b�)�>w�g�^-E&��e�����
�"�{�
��Fp�L�ٺ��@p�كi���*����"�`*���]�X�`����}U4p��"�p�qQ�W'z��j�rȄ���q����bݓ�d�څ���x��z�����1I;���nr��H<4��($��H�hV|��oCg;̺�����>ɗ�a)2b"-c�k���뱌��m͊O�=�|���\�S��x�
�aœ��Pc\a|�߆��|�7���Q���Y��I)G�Y����Y�Vc�S�&ʂ�ڶe&sV.���s2ŋ;ng�!�1Dcݿ/pSqq�/�4p*8�e�o�?5U�*�̇\z��%z�Jӽ��9Y�(�=%n����8K0���)�L.� ����+y��f?#e>�J£��y4�PW�e��3zq�H2a��+�H�I٩O³=�!y28�u�"�YI��#�� ���� Y2���U��Y�1�d��r�V6��A�IUa��Qyq�C���&�HϹ��F>����f�oF�e$E�<U�͟@\�ɹ���I�]����YO۠� ����i����{�r����W��������`�S����_{ҝ<�0ΦK���]�,�"��/�	��\���+���`�;�r2=��#ܤ�����hܐ���87ͦK����s����u���6�"ʻ�cvL���뾬 ;�_�ex��Q�l��Oz�X뻄2tڶ��[m[�Ţ��qWOmL��P�ީ���z����(_�sY�2�fR{�أ�n|5�L�x��x:z}�����1��/N�j<E��?�aV�-c�'�S���}(�]�<^�
���a �
9a�L����u������� M��z��ȼ>ͅ>J�r�K:&	��˸�'�@�@ŷ�����C��L�r��©��A�3����T]f9�Q�kF�y?�����i^�8�湌�ocD�,=�_�v�_�х��'a�MG��ԧ&��Id5�&2?�Y'ݲ� �Z	~L�5�Vi���������7́�݀�����[
�\��]g�[�wV�fVp�Z�V<>䈘N4����e �ڰ�w�(���V�堇	���Nk>��w����e��R�4�۱��mk���GXB�bo�x{Fp�TJ2�m]�m'��U��ǯWTP��*EBaȅ([��Ot��a�3]��D��E4����~h`�!����F�t#��}d?Nһ�jX��-���,��	�*�4�}������0�{U�G4"KB�@�;(@e[�S[p�T��L*�'���?��Aȹ�UcK߁���G^x�k���I<F%ݹ��5Y���]���$�D�Tq�h��^c��W�#X0��s⢒�!��\���i��9@�P���6@<WY�ޱŔ4B �y��g�0��0q�}��f� �܌c������s6Ӕ+M�*���e;������.�w7�ق%�9����������_
����PQ�8���r���O3�H߾���<\��X�퉊f�@
����rO��9͖��W.�.��؛#;������y�����,$̼�����CoKnfȲ
��k��^�/@�`B��D��cTH�����D�'��^~��	E�o�����D��.2�+5^��'W5	���!������[�V>�%Zt�Mu��o���M&*E�ӧ��p�E��F�'�`�V���mJ �%� w�w��SϋL\ְ��q�Ԭ���W~�i���JY��+x*�;���Vꟾ��rs�!�ٞyo}��FJ����<f9�Z1��ǎ��w��=��4g��������]uB[AO[+��7�I! )T�I���̋�YdġF��c�q4�y�>ZI�^�T���|y��p4�1ޥ7��\��+l�^e������q��n�Ô܉@�V�6��XjxI�Ķ}!m`��,X)]:7�6��hP�h,�[ͤ��c���q��uO���`*v=y�
�t�b(B�����ȥ�D����n�4�m�F�~I~ãKD�����N���R��f������P�Q�Է��9����^02I�td�LE��o3U�3+(%�������/I��3�-��0�T�ܫ!���,���P������L>	{�A��K�=Fr� Ξ([W�j���rs��:�ΰ��xZ�D�V��&H$x�v��MU^}D�H������sԱ��S��J۴�
��!��u)��"�B�C�y*��%�Z^-����(�>��|]=���)�S��h�� N5��f�&�9���<����-���6�*�/�e'��Ӕ���	�xz�͌�\	��5�\B-]K���rzZV�`�-7�m]�X�=�}օ.u[jЉ�T �����Sa-hZ>f�T�
������5���!�1I��Iqi��	Lh:�����^��m�fز:���N8;�� ~F[O�	B�N�y)����v�PZ�J��UrF�$P##$8�|��[�)d� �aebکm�4�9�:s���G��`�g��H�J,wX��;<�^��NY���{~�?Bu���K�F%!2��do����?Sn��F9��W�\l�*�#@#�3O�h��'yW|���8�P1O
�KePQ��g����;?����h��W�f�IZujij;E}�`M���3����:������	��L��S�68��Р�4E3Uw4',���_��	�c���~7cz�r|�C±֟G+����i���T�j$Fl�i;�e	�1DiND�O�g,P+��S������ҩx�4@�{%F�u�$�f;7�����$����Y��R>�5zeN����1�]Gy��+D�N2ЏV3��<�_�Z�
ZVO]cN���c:�J���bU��_R���	f�*�����}��伉?�Ԡ�;�N�p��3�k����|Ё�$����a�L�=~�Yl	���l䠠�1���'�NT��xC#�!�����9�2��._m�y�	L�oܓ�����nj�EB|�~Lop28�C9�Y���u|#d��'�1_��U�Ukyq��nb~g�CosA&�(p[����譑m ��0�V`�©d}׸*��� ��ϋ6p��1�K6n��.������:[�b`�`o��ΞD�Q�����ӫDF_%O`v�h�!t��LWh7��~��g����y����>�/9\8�t��l@7t��G:C5�ZG̹9|����C�܈����U�峟�t�5E"ј�1:[?����RJr��B���h�4�<5M<�H��_����D�0Ԝ��[����YZ3 @��U_ޣ�q����!T#�qM~���õ�2�ho�0Y�:��F��X/�-��ѭTF�G�F�!�2 �.�N־�# .�~*��}���g�-Y�-�VnVO�����mx>~�l����Q�gc��ASF�4����PҋV��L�|w�S��g�^�\�l~�b�4Pwb��@���昉��>��]nwV?(}�%x|������ۺ*J�/��(Y,�(�Z)�2K�������K�CPCpa]��E������/6d�F9��h���׉v0h޼�@}�xǶn�yޯ[�
��Z��W�,1S1N��*� @�r��"wjr�n�D�9oG�w
�2�C�����Bf�s�
��O�������[S���̞R�$���G~������$5J �Y"��'	3��m] uV��q8: � 0QTGEҙ��lT��H�.�m�5A�J�C����'�I)�v�(�LEA�0�JA��ٙ2��]Cq�yyғH�4'�'����ѐB	��}��$>4�ٜ1��B-a�;҃����0��B�a���ou�W��S,(�&�`C#.i7+M�^��|�%4t�3Yu�|�!Mi��Ow����q��q�`��u�"k��_d?+�[�\�g{^oU���{�>�݈�:����f���]Cz�����:�Q�]T���U* �!����yl��Y}k)�K���,�#0�Q%!�V�M��9�<3zv�ӕG[�)��:���ۓWϸ��7��
?�ͬ>���t�F�3�sR� �P�B��z���l����]W��F��b�"�>�1�=���y��,�k�Ѐ���(�B���	|�{D�U�s��Xȶ��5�t����0�\ܰ���'؉���r��)�Da0��/ML�x�J�yܑlپ�9�����p�Z��(�!���ѣ;Sz��v9?@��WQ�V@�F�E0Bq�(� �� �z���j.b����H��o�����Z���:86�y?u�N谹[s��)!����ˍ@g�N�COQ���Л���K߰�-]�ƴ."PVg^j��^̳�q(��4��|r��	43�2{�F�˳mwGYl^���Z�0?�� �&`ۿ���~�;T����!l2iljKF���6����ݚ��9�y��'x]]�Y��Df�&�/���*]�+��)v�Z�H+��؆���= �,K6�M������%���qh:�5��H�����y7E���Hb=������I�jz&i閌'��� T+v���;兺��۶�"�6f�f��;[o����6!z%�C@���,�5��������6G�01�MH���.����(6j�Ȝ���n{%&���_�<�q�0��FZ7�&H��)�)���g���"��Fxd9��mQ��(��Ϥ�c������n��=YT? ��~��a���׫ӎq+�21�*s��NP��Z(,����O�����&^��l<?�jC&��MQ�0����;q���+lE���c���mu���4�G����1r�����܁����b���6��9}����~�X��x��"D�s�=���]�To|�\�ZjeAjv��^`o��:r���pk���;��hG�Uui扩<-��u,8��[�  �s`�D_�8���f�w&@@���f'&���Oa�j�N0βk�m�R�>q��u�Ψ;��X"D�&k]��Q�7=i�A�ɹ!
.�q���װ=��)��></�����'�;^l6��~�&�߈�vYu?ڟ��/K ��@7�#fO�T�$d�ݚ��AתD�hzGp$`[L���^�Ø�n�� =��`S�^�T��7:�/U�ߌ���A�c �E��qY���6���'T�)�Y��bzЫ�hA�<]�a�i�"���5YF��Z��P�\��\��v�\a&�<Q��Tn2��d)}1$����s�S.���]���f��ngC:Z��rK� Qͺ �ah� t������������E�n�wi;R�����w�8y����+i�ˈ_DDpq�7�G�Bi�B�u�IF��{��d`�������tT9"��M��vt��;�]i�G�]�N��0�&e=9�b)�߯��>��(vT��K��ظ����q;�A���7m�9z�_��;&���ѕE�LI���;*�qH�����@�IB5�j�ثCl��Uɪ��V��E|+V�C�u�B��]گ�1#`mr;،uu���ĕ�����5}�����򱽘Ԓ�X2U����=����
��V��0���8%��[��Vxl�hN�=�l������=�\��	X��d�_�'��Il�����뢾c`�9�S�o�׸���ӯ�컓 ����E��"X��G�c�L��M��6�#�������ӡZ{JwcM�2-}�=m�n�$����5�T� ����L���ND��Ԝv\Cy����S��w����yE�Q5����7�I_pO-�m�fjW�>W�"{��9vV$�]����]>4�u��{��0�N��h+���(J���ȥ�ݟ������(��`n]����K��9�C��ߤ�6c�����ʃ?B�:}̀T���g`�w��|� Pj�$>D9���{Ay�G�d�?���*��q#�[��VB3* ���a���:�џ��$��Z��P��KN��=�p��3h`a��`���ux�$�)Wg�ˍ:#՝"���w���}idݼ�5"H/P�f����*�E1�
4+\x ���p�*8�����_xF����+��Y����NW)d���%�-g��ZwpG�/�`��p%i��0=����*?�h��=�n���A_.O1�,�ԗH�(C���~-Ј�	�Q� M�NgX\�������J9'�т��nV����$J�T,y����e(@ޝX���O���3�Q����Ue�n�m�?D>P�4���Ƶ��Q��6&��Q���J}'~��#)���R;�e��w0�l��즓
pagʷ���E>{�,t��'m8"��.j� �6�yM@�<�}}#��F見��~xh���jŔoH4i��e͎{�H0��l�#���Co���kќ9�z����s�n>"�ɰ�v�iR�m5��J��%y�M�HN��+�*���ۨ��[ă �+&|��T��\���M4���STn�VH
�
%LZH5VwO�P_O20��(y��"^�Bf2�nP�t�\G4;t�� 6��hՖ��}�����r��-�l��sWn��A�W�*E2�o�	����j.m��3���W�k+Jس��	S��&�*����.���d	�姸��.���J�aٰ��r`��6=q����mz&1��4�Di6�{[��ކ��ߔ�f>��H���*�6m�@/%�5�Un�f�m:5Ɂ.�1@fΡ��T�G�?f��� y]o��?X4晤����e>��ڌ�~�)*��� �����eCO��[%� 1�>�H�_\tچ*����%����MM��?����K¹���_p��[y! >�$%���v���3�?:����� k#{�JL6���P�i%�U��
�F�0$1�HK�-�Hj�&OZy`P��e1�jc�/D����c�,Q�DK̀B��2��'^u+f:�ei��IFk���pL�#Z��J,\|���~X��	���M��uup�����a��mG�����Y��b������)j�x���Z�E_U��-O��,�x�Q¸Zޕ	��24Q&1O$�W��,߉���r�B|1��h������[9�����!�sL e�h��%FZ��n��s�Z �.�B�^*��!�]Ml��(���;K�al�x���&���|����ﭱ�n�����hi���,���HMb�n�:[���KQ!� B��}����
s`Hy��º��l��?a��H& M5YL�'K��}�Yi�y>����sk�LGE��o5�u}B�S�ax�M1�iF=zW`k�)6����eG�p�R�5���ֵ�<Q�|�q�Q]ۑ{�a��&s>s�!!0�uT�b��=G���w\#:!�qM���ٓ�C����NMl`E��PGv�^E��h��zQ�;qA����<�6~��x� ��'8����D��b��)���۔tG���G��_9� �+������7�
!�d$<Wr+����Lx�pb6��R�e���DDEh?��5����]�!>�l5?̶/����V��䍳/�=��K�̂�Xs!}�]��#Tܦmg�20�V���Ѵ�g�n`�4[�</GJ�u����sCz�CKaa�<���)oRn��h��S��
���K�!�J�ԫ����h^�pZ�6��X������ws%�(Z	b����W�啂��;$+V��y#���|6��C"&��3�-�-�����8����엝J���ּA�'��-<�u_%T��%"����d!�m�PG�k��}ꍴ
|yj�[� �/����4d���܋�gG�A6����uE�7'Ԩ�nm��v��5��Y��D�31|�#N��0�vǑ��oWbVG��M��[��JL��ԛhY�]v���/%�� uҮ����y��
���TuHx��zZ�,.h;5p���(L�5�j�>�Ǖ���L[4V���*=4a�y��I��������ja`]��� cIc�9���i���N�Y��ħ�=dUm_�ų����2'�/J�$�)��^|�W�EI-$��惛���f�(8�=&�=��ó��5zM&��<g��0��I5��gb!�9W\�I]��Y���x�/
Ú�[̛�@lm���9k��j����Ȼ�7@,��|���E����9�?��V�=��K�X-�w��F4R�Հ�;C�J�J�ro�+�:{	T���l�<�5NB�@{��K.�{��-TU���;�.���Op�G��H��`�x9���!�qm���g�V�!���������3���ݙ�/��>���?�˙�5�&�y�Z�ԃL[ꛀݵW���Y�'Rx��HP�o{�:�	�2 �*z�	��t9�<  ]\����*b+8�u� ʭ	bLG����m6�3��|��ğr߫�� ??=��.�O}b|���m����Zoxꐸ�bl|�o�Hk+���s�6�"�i�MC���d.�h�<��1�g$���N}����O�Y�l/Q�4?�/��
(��^�j�����������جc"7m�A���L�2H!o��?�+��� \��0�5rA�����;�2\O���	s������������Q�Gyߙ�+Щ"G��6%8�7{�Y����4��g��oٰ�z��޶W��=�8����
�? $�+�>C$���*��}a!{߿����-���#ǕDFcy��N�3�]�	_U��Bk� 7�}{4_���4�~ c���n�̭�����V&���F�&�E("�@|�:86M��ι�,�f�h�;jf����{D�5ɔ��:3w���A%�(nF%q�y�AVzs�6eB�����qJf��=u|dadY��dv�؎�pn&)��[��\�l�����!��lʣ�u�K����ח_��EAn?�U�Ҹ�g�2:y�!WP�y d�4�[0�N�8���!�� ����3��.��&��d����e���a��|o�anb]�^\J��w��V� �ݽ�b+ό��ro��/�l����b�=k��g���	80*5K$��zn]`�sW�Z|�w�eʽ0����f�A���0j�,�ZF�Ͳ�N׻�E�5�h[,�-AL��� �_�	��"6'�G����]�7�Q�:"�8>�x2A�e��-�8q�̓��Ш���d��`� :k���/��{�h�Gh�g9�QE���&ڨ���_����ƣt���y��D�@T���"L�=��nL��O�l3���:�mLl�2�7�U��ńw��'�L����Ñ�T��
��˩�Z��]�}t��vŸ��0�2�z���O$o�4F��Q���Ru�;0�՟��dW|�<
h	9hV��)��i��\�M�����
9��g1
���"�[ϗ��O�Z{�[`� �>�i����jWqF����n��M�|�[Br�vY�D.T�>��6Gg؝�W7i*�Ìͽ5�sY�Z�ijdBQ�
ea���lD�D)���+Tv4	��z�&a�0]������Ǉ�*X�}�Y��,5 #����P��-��"
�2��͍K�U�}��� _#UW��o��Ѡ.+Wv�U���ä:a2�Ѳ!���	з�t��B�5\-͇ύu]2��ȦK��sR�O/�ʞp(]��i��T�!ı.���	�qǫ�3�/������Z��xO�*�2:�
PY��Z��ˈc�i��:0�w�0���v�l��)A��ƻ
�6b��9��J���SD^�N��T�=E�{��T�{�Ch�� d�8�Jc�`�װ� *����wl���s��3���^g���;����x ��^TT$7\����6�>��b�.��+|
�3"(�c+�g��[���*1w�f7�-h����Ĭ� Xi����(#�Z9`<[k%p)��}8O���=ߵJ4t����n�cf��tc�!�,S�a�ͷz�EQQ����'�c����uh��a����b�蝧�R��X����$��饋��*��F9~A�,�z��~�&$g�G�"Z�k�˵>z��#���j�iU%lz�K�WDv�����!=�t�<���;F�l��;��/i���J'�JS��1���K��]�榦�,@�C���FS�y�V���űE���]�%RN��&�Z��'�97��W��P�ޙ���y��3�B�6L?,��\��-�ny;�ш����Ÿ���'�+Ȏ˰��?��=�'���کWVl��_���B,�FY���[��Ec*�>�O��n���1�;����y��~���߱)@1mb��Z�f<m��Ӊh�����.�ΪW�����٧�X9�RT��b����CM9�tJ��u���~�,���v�IaB�I0j��eG�Z���;4�0k���A�6��u5�ź0�T�,&���-��!�ZmP�c<�3�r%�/<k��֔/(����������_��(*�Z+``�#�-CD6�����}�.��t,�X���Z�����
����'��#6�<�
��X�I�x߉�4�-y??>l
c��kqˈ���ѹT��ū�bOXD7�b8�KV���'Ad^��2�% |�a,a54aX��Ӎ�a-�jt��"H�*��(��,�|�[��.>|>S�/1���G�%��Q�d�4)jk�@���gy;�WqV��m�;{�Y��|Ө5z��l��jZ޲��� @�D6�*�p�3�#�A&�E2�)�!xq�K��S�s�,�ᓣ(���&���h�P�{���	���GL�=1�N�B��q6c�������\��K�>����h^�e7����L�W1���-\���o���.eg���\]�9����Z˓�tm�i ��m�p�w��G˾�|�RoU�5�ܨ�����v�ɶ0e4����Z��F��}�HP�6���~��E�0�z��qTey0�1�4�$��ޕ��xeE��j·E���,5:�?��*�����(�ܘ��Z�9f�jF�:��X鈛t�I�'�j�K2�ahE�w�m	
f�ĝߟ��w��/VJ��ܖ�~����n����+���Jp�wv'�g�� Z�L��������F�T�$�)������K#>�.w��b?��]V�,J�[S׃��&8u��e�
*�i5�԰�!#��o�N����|oP� ����Mer^h���Ύ.1�95o�P��!z d����-��źy'D�)��pݎd$����X�V;9�������8&�Q�u�<��ϳ�j`}��6�m���?I��m�� D�:�پ�E֠gD��T��e�:�C���ms�Z���
����e����e!:B׶��>qhw���_�(#�c���?���h�W�br�t��Q�s!?�t_MD��@fs1�C$֓�3p�-����t��ؖt"�����8�,_ӊ`��ƫ�<���)�Q�"
�̹��7���p>�tp�TKɁ�������a2��Tih�iKO#��H��a<�k(\~x6q�B�1JB$S�g�y�r�;��h�b��mf�v���o�_�Iw��"�(� �H
Ro�-c%oI��|/��l���:w�&o���9������GV<.�f��ܓ_qܽ�O��6�xvΓ�f�?<��4��֒y*^_jM4�#(��f7���\-�ؼ��r�NvC� q'��h��\xL�O��Li�*-���w�+𑰚r���x;��'�Q��r3��>��&3����B����e���ӭ�EF�����(<}e��r�{�
�Z�8Ji���&oE���gz�>��<�fXE?T^��a)[�!�U�F���o�鿷�k����b���0>]�R՘8�m	Szڮ����u(~p�r��eӺ�3��I�_6ߚ�
�4���Fܺ�@`ypb�16�n~qG"�e������A�����~��c?j iY�EC�O��o�]rM�✄AGF��[#��[����ݕ�Ag��.�vB%,�S�b�A�ҥ��ǪT��(v�9�AU���Cd�H1�~��ȯmӌc�թ�̇�b;��F����i���=�£�W`_ˢ�J��3qr�)�)B���U6�b��z~��($ up�V��A�S��¹��xǪE7����Q�h�!���u18�&w����Ń�_�5�8��F�09.�Xܼ���ɨҎ��Cc��h@���5�����Ɉ���N��F���}L�&�js2>����/N�S� ��޵���<����n@^�*iccj�B)��Mo���_c_3Γ�3�m"&.�JFWwY�����!���B������T����ؑI^�ZH-�:�q<A��p�����@ե�W4=^��g~t���%�6�>�Ҋ,�q.J��|��{	=Z��;rMf-�)0���
��@bE�p�T~�t��a�AE�{��[����.�iՊg�eGu��S�!�#qD�g��6W>�0O8y���$��c���W�3��=n�\�CƮͰ��Й���s9,va{���w	e#$b�/�1�/��s���3R�qu�[n�����OT���4�	7�6��vS���Hݸ	�D�Sq�5���K])Z��Ǟt�E�A`I.FaʓG���dd��g�bAU�XZO�������+��YQ<R��q�����%���!����8#��`������O8H��3]��`:��(�wi�R-I̅m��^q����-�r� ���_c�1U������8�{Sk�wf��)�u"��Ǆ�6HdD�g͋�R�<T�L&�uYϫ�I�� դ#��<��q_n���j��y�b������$��l�%����!_��z�B>�^�f�#iOmp-l�YZ��k�@��y?��z_^c�VØ�{'ō�����WjUjZ�o�┫�ct
E�
#���8i���y㒬���:&I%�C�C�a���G���*ߣ���j�c����/�n	�5y/�{Q�b�����-��\"�F���P���;
��T�`|�/�\��"�>I��`�z�4�- ~�S�F���C!XA�)l0踊x�����>���h@ױ2)���9�|b��-��"
��V�����^@��������"?�K*213�w����`I���y��*�paNC��%�͓��t�=*�� S�T��������˻I3yaXCxx��%5��ȇ��-�L	b"��&��^�Ά�k��:T��	�j�E*ً�-�׭ƿ&�m�Uz@��U6h�Q{������k�������pyCβ]�����ǫ�f�?�<�?f4����� �J�WJ��מ2�DL*@�!���LIJ�Y��M�2�&;���wg%��ON���x(߂B�r�l=��^1]��]v�8[�V`�G���xZ�c��FNmJi˖r�Gc�g�t �L�MpA\�q�3�q�`�2~eH����g��� �P��V�V�+����t׽�msa+:�u���_�x��yr/�h��,��b����j6 L(n��oI��xe�5C���n�A�n�i��#�5T�.���[	馾�_��)!�IbXvxEH�`C��������+�	y��P
*\�+�9���5(=�x�~��d݋�:6EUR�V~�����iM02�/B?L�9c�u��DH�X���������������NUN���\��M<Z��=xT�Cm�VHR^� �P���th�+���FzI�%0���?�	�Q�qNY6O��`sr�����H	���*9}�
^B�Uvj�ah��xAHu��Z7\4rO��7E���^m���Դ���cK��`��G�ǥ�l$q-P�X=���ak	���ɇ�?#���kK!L�h~?p�+|�_�_V1�y�!�zW��+p��f���*�ä�^*�e%�i��خ��|�m"in�����}�AuO'���(����Y��mU������ff!}p����m��=���3�O<ݒ��B *6؍*�m`gκ�u͚azK�'̴͜��.��Ub.��/]<E\|$��CP�0�ծ�P�e����u1�H'�#	VJeoo�=L�ǯB�r�s�!�S_�ꢻ�:N��'z��0�)>H�Dݻ��7�؞��˻�Z�KY���"�2�ڞ=��~��9jB�ҨB^l����=���^�Ɏ�S�:n�뚊�q��4��B���@Y�u�Y���/�1!�%GL��M��HeJ�M<��� �mæ�������cWVeQ����N����G�N̎��v8�wCT����ݯ������[�h�/�Ǽ<�;�g�D`����A1��@�2�^�����^֞�q�WU�YPh�ml�w�Z�Z.�j>���6��$j�w*8�JgE��g���q�A$��z�C㕏�<3z�/��lm� �O3`�+y��s�p8{��_o#VBU:SVOp.�O�s�*e�B6����tk��ǫZ�\�$3�[��	;YG�ؙ����42�˻<N�����}��_��ݾ�C� ��4xe�j�R�$�.��?�iC�.y�k=/� _�@��z�pp�rP��i�m�r�;�R�?���>ԩ����>aIIOf��p֝D<��D!�(2|��dƕ���B�Z�����i-{�;���d�g�&���u�q:�F×��>��@P���u��$O-�����f�)�O��tn��#�����=+�&x�@FQN��-�	F.^}���$r �V�U~�1ϱh�����D�"��VD���pC�"�����F����h�wbt=N�l�M�q��Mq0p -Gve������}�q&UD���;�~�|`_�w�׏
 �뚰������)&TJO=胱��}���ҞdW���%���V���,i9V�K|��T��l�Y��٩�i�	�֔�`|�	� q�d�H"GV�$�|�M���z�n�;�xɫ��V����G!��G�&�XA��r�S�(q�o/$�ד7<|%�E���ɡR�b<�8ـ����l�_K���"�5&��cHN8�ucK����k�Ov��R�F� >^�d���k�l�XtǓ,h���(��u��u�����c?�}D~�����J%-|Q��RF�)��`E�/�mi���<�
�©�$?�H�� �OB���R&:���q�]��
�e��x8�|5���󘻐��@}��o'�җ��V�-my�$�z/TQ~���Q��L����4�$sJ4/)�Jj`��BAQT�07������e��������]��*���P?��O��X,֋�D�3&t�乹r\����v�6$X�R3���=g-��2��.��(��&b�9}�[F�|ʢg'�$	��B�e�����D�#ѕ�(%��q7�
����Þ��&����;��j���} �-���,S懛��E<����?&I6w�V���Nƹ����q�L�$*w���������c9ď��3���H6-O�n.��Mچ
%l��an����"xE��}��6U�)����?}�*�R�[֩{[iQ�F�BOM-'��G�F?�M[8&.���i567La��΅��t�zmc�����ݾ�������Ц������;�7I=�4���2EPRa�g��h�~�J��󜡾s?;���p�Ec��7����k]zX�;��HcFckV�p9�-�KE�n4����A�?��ݕ�N����<��$��1��cx�\�Y.Ʉj�ۑ$EGk�ϑ��4�����,���(�7454&�l�扤�`��t3�^	<�uI��y�/��b�(��fS".��/��d�\�ns�D_ ���"�t�m�(i#6�
U�Z"����x���W�}+��{zsr|����c�SC�����v �8���R�VD7�L�7�s �\ ���ķ����EcC��܌���"������sdyrWa0��0*��0�@�\�΍iW,�����i�}� �hwH4o�]�E[ ��=gҚqw���G2��#���bg���en(�ܺ�:��4Z'�V;�+���5����M��U��AU!-�#�%��ABZq4���\T���D�B�#%s3X�>�ab)[`T���]��]���D��'��4�N�k����sV���TlCӝ���:H��8y%��>=�p[:Y�Gn�ɉ�qۭ ��TV�q��JсT�U�C��ʰɼ�YA	�@�z=��K�&J�/v�'��� �uyiD�ӈ3Ex�u'L����Є���P��T��΀���b�
��QM�B���U6.��i9�Qx�Y[���M��tɶR�8ѭ��9v�9�`7�t#�C{��9�y��%Aj¡�����\�?f�sp���G+O�D���-C�ܞ�!(Z.F,/7�d~�&�ϺFe˛��6��J�M��x\E�#��<�/��z4$��]�S�s�%ͰD֔����w�3N���J&̛&�?�yϵy���������[]JzX��
��jF�d��!�Ⱦ`#�5S�B��F��� ǈ��C�!YB4����]R��Ǳ�-��L�'�;�s$a���˴ �����3c��I�P�5�[�mt#���;��s^H{D��N�cB��Ù��\����&�r ��U7ޒ$�T�@��kS���'�%́���0����D�쪔���j��|cM4���z�E�r.��p'����$��=9	��qS��T�z=i���>���MG�q��ڣ/���ὺ�AǚSVV�m���(fA�k�l��WΜtn�#��j9��/���/���\�d;��O�o���>�[+X���XדmU�v��.��
=-S{�
�%�(����� ��5Oe��R��W{����>L� W-�b<�
��� Q61�zO��l:O�ԚMT',4�b��E��j�_��``Jڎ^"��u�x
ǅeU�0�!̔����Y�Tj�� $�h�>�|�U�R+��-u9�`3��P�D�d�4��$Q��t�����Ġ�1�ŶL�jT�ys����ɦ��>�%��y�#R`+���d]����#_��#O�S�N4[=i}��e��jA��a��o�"�F|��'�'�����_Ĥq޿Kjz^1�G�H�H3�#��3@�uU5wo���j�G�W9[�ؘ�{U�2ݯ���m�_��Y��D�Fkd�	�Ee*<M6a8p��'��Z��'L�(�i�iO�[�2z�$�#y��n����*o����g!��~ҾQd'd�k��k�U�&��G�:���e͏?���uQty
u�%Q�.V�I|���[��h]w�Lji"�z}[ơ�h}��?�P�|%�"�6�3��­н�6h�\a����9K̅l�^����G��tG��h�e;�B�#��i�5Mr}l�/xh��!F#d �a�1܃3w��\;��)�#�k���^�o������׀��,f(Ʈx��.ʈP?�_��$4��{<��71�٠`���m�)ذ�d
����TeO�߿ $f������%y�Q�(9D�}�݊Vv�왌�CZ��>���I:H8t_��H�kѭ��n�s��JdR)ikq�_N�!�/��'�o���f��B�y�HH6�t_��O0�q�Ǜ(��g��]��i�%V�q3A�{\��c�
�'�xٝCJ�灜"`\�C�`�x�`J���vP��9���P�*�`�)
�?���5cB�)<(�C�����u�
�qoHp�N�W}�e���#71T��J�Q��i#�.[2�:���<��Ffe����Yh�d�S���F�$�X���o��TOfu��������4��6��Q�`���߹�q���ۛN�\f'x��=X���MՔsO$�d��-�2 ��Z�ր}�S��c�4�
"�w�f�n��P6�~�#y��HlN�ET~���k����#o����Vއb!��j��f:[�U_f�;��i��KG�9 :�IЀߕ��B(���Pf��~�F�HwMz��p4'�KA�߮�Z��A�ݱ�*���k�G�~Ux�h��7��w4%6�~ҙ���6�w����lj�]ώ��;�ϛWE[S���v�T����@L��s���me�	���V�e��b�j7�W,V����'�e�1�[qm�G���Y���>�n~��׆ra�.3氭
j�4���VᆼMA��O��N�j�����.C��*�����#��΀�bn�ఖ��L��X9фA�Q�k�� � ��N�W��:���[މ�D�6� �ἂ��1����U}H'V��B����p����:WoGk�	.�_�$d ��árXh����j��4��@�؀�?�3�ҁ���Y��b�e��#�4fwh0�C)g��~>��}.dL��E�矎}�" G�\�Ih<w�D�18�I��bq�
91�H��Y�� ����9�%���ƻ�3�f��'DI;�km��[i�O����B�52w�m=�B�?���()ˏ���܂^iRG�k���b�DKβ�H����Vu	�zNcJňƫ���:�F������>���-����r� ��s}5W�
�ˤ�xW�� ���s"�p���@�^~�8e(��k���m�޾w�����b��F,/\1�5�����о�ñ���2x3��	og�e��g�8�3Z�J���Lt��k���<% 2*���,��U��%*�{yw���/jZ�ޥ�oj�6������c���X|

���MR8.�"UZ�N�4}�H9V�W�p0Q}��ǞK������IFXPI�-Y��x�^;��I��C����؁�~�'ռ�.����1��^�`1v?�ɤٹc���+d���ʎ�JH{[��Øt�ݵ�6u�<��e���U�}����I�#�ŋs���@uE�#&��R^��4g�ꥎ���ѐ���bQ|�;��
�uj��4���m5���bxt�ȧ�D[@��<z����x�ML$Q�ZH�tzfҢ�/ �����W�<�Az=���8a6U?"�re5Ȅ,����	W�t�[���n��J���dӕ^v��n�ę�_,�@8�C}	z�Y��#�,ǍZ���R��_T�۷��K�(����)�S{2$�*�4�D/LLWC2�H(Ǔ{4�K��޾!Z�ݣ&�q=˻v;�m�sL&�"�q�gR�l�%6�����0�@|Nz�a1m��E��	M߯���(�q�����?c$-�A�^
�Fί�ѣf��IX� ��/sGw#�X;�b�l�=u�PU
{�khgϵ�g���߻sV����gYƏ���'��t���{`qIb��7��+���B3��ݟ��'nM���9��J0N�$�P�%J�����4B�qݻt�1zaF���$�̾y Ʉyi��5`��:�K6�`�����ߊ{+N��t!+�����{�b
�͌����!)�X�p���|�_Հ��-.����_J�:�m��o�o5	ASl�xH@�IflG{�*��:�l��i[M�{鷕�h�K��>2��z��f�9��?doI�>�G��׽����Գ����rv���&e��8Z�OLM����Ȟ-M�^I��6	W�R���8�J�=����x��2��"�Z߻��鑽Ϗު�C��fUc�+/V�3����L�*7���˹5n�����_������"�_CŮiiL~��O!��Pi�Ugy|�vN0>!�08t$��l�:���� "+6"�J;u	��.�c�'0g9 �e�y=�h��Y�c�wv
�����K��	*oM2rm��zQ�8�h��6%����݆�,c2�B�ذY�}ϸa�~I��z�z� o���^i���ŉh�����!'��HH�h�*2#���'*�5�Lk��SeP\�7|�!Z��*�[>�'Y�-l���f�o�:��΅���=���=R��-��1�h<<�"�`oOVc��4�R��i{�8�9S�#Ҡ���܎}���N�:��]K�<���O��b�w,��d~{�i}�t�j��"�멉<���l��N�]������Z��}����>!Y74�W�LŅ�Kک'\�	i�(�a-NC��1�zS���I�kG���a�	>zofZ ��z�|~����6b�
>�������e9P ���+�dġu>�Z�<�`ZS(��b�����
�ȚV�ؘ��i���M�x���)4��֪��,�+�vB�)���N����=4�`���s�7S��~�-Ϲ"*�%� ����ћ^��?������g� ���Q���kh��ݹ��{��S�OU1$��4�2�]K�EB��׋hlT�Kt��"���03¬DPN��W��SYއ� w}�bE�ᐰ���`��S�1;]E;�J@X�B���8m�кY?�X�+�6Ji����EZs�r�xw���A�T�0�-P���B�Yts�>V��,�U�-�I�T�#!�����'�}�Զ[��)I5�!Zs� D���)��Ĳ詨��
m�f re3���n���ߘ��T�rQg�K��,^���>�wjM!5���2��p2�j�w���Iw-lВv���dۤ�!��������f�?&�Hi,NOJ�&�����;����=#�!���5��LȏiH��0S�y��T��V��M?vW<�&r}����{��D�)*�󇐖�L�|_b^��K���Fa�����G�6��n�d���e�˂�U��1_5��8���	޹�|�vo,\K�����s:�GW�1fi�}��i&�ܳ��ꕲ�i���i>�Th���QZ��j#����,�t�L��I�e��Ԕ����|�2/���箦!��R3���үV�RP�4{�s����?�͝>/�M&
�����{H�\*F�G3#��gܼ ��h���3��if�_\�T�	ʺB��|����L�m:��s�U�-,\|�2MQ���(�V���@���xPz���D�W����i���k~�-�s#�����Rj/�F,8�lF�=��r� �^�ʑ6���V�.�o%n���t�С����HT�rjF�^;�ƶl�J:�Z�]P����A�&EWp�z�>��8�5��YG��ӷr��������Z�,��4��TJ�k�4���TzL֗6	���Z4����R=o�\����� �i��{߅�{������t��ok̞�ב�Z,���n���� Y�k����g�E�3O�HK�U��F��f����9���[@n]�b�w��C�P٭J�[���0�?C��xƈ;L��:��0�"kx"��6 �?�eb��m��Z�����h�A�	Ἁ��BF��r1Љ�fN��K93J;��h��"��C��C%x�g>�4����k4�T��SF^�Pw,���~Lø,<�{��%*�*V��ބ���bTH	ջ����+W:B1"�^��sOU,��H>Tb#{�6��L�o�Uz�k�D�n��)SC�l����vN�S�y��O�c �s����D��x|�hj��3!\Ǎ�LH��[v�~�s�P6.�T�6d�Z~Q�F)�!ȟ��#*@�m��Jl)ތ5���H	��>�X^�;�7�ԫ��{���s8/��*Y�PB9���������
d�*f�"��
4ҡ/{,&$s��
�e<��ho$�e�j�Q}_З��J�հ��X~��F�e�W�<4����>Sj�����|.m��f&X��i�g�n/nY�j�1�$BO��s��{Ҝ��	P��ݨ��c_�ݣ3z�`z��7}1�.��6�]̀M�q�ay��Z�Es9(��8�S���ռL���SO�ku(�]�z�-���S�����t���'\�zK|t���eU[�oK�����yJ�<�Z­	Fz-qD���ߦ4Ǵc�|X]�Hie8��uy���j��Foɀ#'}D�v�@1}��Mд��m�8�$b!�*���2I(���sfɎR(�='A���@����-�H�H�CZ�)M�� qt�U�K�5�ѕ������,�D�����b���kAx��K4LF>�oc^-�T %�ov����N2��-.�����O޻]j�z�j
���4�4��]�@Q�Zp��͗-l�m����f�H���j6�D�����n���#l6�ȭ���A�����O����������|%vM@����g�)?Gs�I>�9Óٴ��1挗m�T =g2+��Fuf*��\��Xm0������ J���d���K��(�����:�����ɒlbs|�<#X�ǒ�Ao}�f�#X���g�@ܐڝ�Pm�8��rgg&ԋ�P��V���~#A1YBd�A��J���7-S��>~��E�k`a�:�t����a5��)�˲������rrj�E7fc=�ņ ����8X��f),�{T��y� I�Q@[- aqm!w�NU�{{��,�B��v�/�i�#m"���G�Eڠ���)�Es.�%� 1�;k���v=�ړ�PUz�Np�3�-�m�*�ޟ���0z�@8�ΈǛ��<L��c���'�#3��L)��S��BյN��K�?V�Z����QK�m�ŀ^
���8�c�f������2���<�u��z��uE��A��+k��mNF�Dat0����l�;m��I<:����f�(�Cj>��vy�6�Y�{��I"�w`�Fzj���zu���3F���o������*�����Lwi��9�F{��b�y���\,����u���Z�<�R��0�ʓ_�Q��[��+j^��#P��61cZ��.�������7���NY�/�'W��d� ��DZu6��On���IE_�m�w���kehCW����ۿ��ü�,��C���-81Z"�AM:�r1�[���f�MK��"���5�t9P��zlp��غ�O;&ef�AJ���Q�����{�^i�q��^v����XDA+��'2�ctn ���d�"�I"�HP�_��4��q�����Q��=��6k�@�qE�#���t6N�7y8����̠����\Qh�T�q{�8���e�V��9��Sxu���t$ ���2���"CAB��gy+2k!Z�Wb/�jL�\iA�W����^�X�N)���+��sRk�<
��\+����r�Xⵙ�ͨ	 �ڱ�������Z)P�_^���5s�pka���f`�	�M����b2ѝ�d�L��[0�����Fvx/~Ȇ���y��]�R�<�|K�$�]�B*[�غ]7��8P�����IɷVM!�Ml��X,�4�a�g-��'ʅ�b��|�+��]鏑�x;o�g�����Tp���%���[7_:���	�z��"�rw2�R�3=��ˤ��N�����"y�TI����&��G<`������1#u���O�F�R�6�����jSV74��w�gj�n7�^z�1+���|�͕_�6��cx-�n�W���I)�9�_�b��_�Wz8q2@[�Y�dU�mF	3li�2;a���)�cyG�҈w��aW�[���L�,�ek��#(�S���.9+�#���Qw�AP�'!s�J���U_�����-���M(��:���ޓo*�c.^ɲ��`��������ы��@��I�)��@�����6=�6#	�e�F)l�wY���C.ZsV�t#1��kp�^Ү������%U21_p�k�~�j���@3LEiZ�}�SYl�O�r���@񭙠�m��C�cEʔ����t�@��(�_��#X��0^P>�s�Ʊ����Tu�m�TX��j%��0~�D��'��"<xz���u� ���v6&���@ �ȏA�4j�h�Z*��<�ڶ��g�i��N @_>�z��Ԉ@*e���!�;�;,-���Y˱Y��Qh<��J�(\8c͗ByZ 摉�_��8�Y�&}W�L��������)��ı���~��F���M���J�IҔ`���4�����E|F�n+>��'i5��o �(�<��\(^��4��OH�=P����̟=���a�J��?T桜�ƺ#{���3I��l�]���8ݫ��	���J���F��i���>�sj/���s���F,��Q@�����]�����	��c@WF�<|)�\�x,�����ZE.B��_�|~ճ�,����/�S��W��5�s��f �e��.>�>b9D�ز�����T�����/�W��&��A�G��C�2w��Y������㍄8G��?\�b-����ʄ���G���+���x�-AF�Яs��3ʾ�?�s�Z����!e�Q��wEHyG��o}��Of҃�Po��Ĭ�4���`$�g�`S�?Z��.�*��`Y,Z�g��fqaR%������4pŕnl�d���$�0:\RCr�5s�4����6���;�T�_��$ƱA{9D\�����&�[��F����X��x�@��xH����qm6��E�z,M�'ވ�2x�K���yO��¤�2��`W���:a�S�ɸ��3�U�`�An ,L�UT݇^��h�<�J�6<e�U��45�3��n�������M����N��k���-�HE$RI��p���\�,��S8p��G��%�Ҫ�*�x]���N;1���Ψ�lWD\3�sΰ���1��a�d��c/�Nj"���]_i�G�܂�S.Bq�1ˑ�k�LcwQ�<�n4%.���Q�kmj��"�b�̴[ ����%���a��t8��7 �ŝ��Ӛ5}��k��>�PZ�&sU1Ě��k3S�ɨY�˅��g� Z)o>:J�@h�,��,}eߔ��N��V�a;m6 �E4�i۽\`RO%qʊ%�&�k��F=���.혁C?���Tk��BI�%�����U=ӑ�I��Ei$VᎹM�֯$�j�'z콈W��jbeHC�6ޏ��}�,L,3L����_ _p6X�]n�*:��k���m5q|вD�})� �I};-o��+�����L4,�>����f��o�	�u+���\�G�@25�PKLY����Lp\1�U� UQ�FUR7�q�P��a>���dz9}i�����������V�{w�����9.#��������⪌�c�_�z�,)-��Y�=��y�5ő�9E����uNtT�7�C6�dX�>(������w��bY3d��`U���'�?�$F���|h��������Dg�@ף Z�ځ���D4�P:�tX��w���_4�	�O�ad�lx��,����uUPǆ�Y,��9����qI��=s�FD�������M9j���ʈ"*%�~�7�a��V^��ߖ"�P���������b�׺C�7b��q~{0�v��� �D�D�Ө�r@��� �52t}�l;X�$�7=<��-�����yh1o�f�vyc���R�}r�Q���{�g���8OdW�8�RJޝ�c��*�]��X�zj�8�h�ar;c���]�Yë��o�ۄ�*�q3�k`$�����6�C=�<`�5�\Z2�$�[�!��s��[���5��+?�P����{�fT!������9��F��g�ܕB��t�����ͩlSkt�7���9B�Ж�jv��:G��P��s�#��r��耈GP�7~d$���9�A1:e �0�g��&����r�>�(���i�{ዡ��x>x4?o��I�{�PÈ~�D�4�hϝX%�l���9q9��wW��,�uH�?�(3(�*:�|h���`�&@*��S��T|���ڀ��2��s��ۧ ��<o	�3�OIt!}��1�b6�b�X(io���?���e種���dq%�v�Me0j.��W���Ɔ�Qn�l�7�B�F-c��1:�9K���� �㫰��R�^�5����dڐc	J��t��xq�d,���``�(�������]&h]�S�_��b���J,���<;��d4B��3��� >��9l���-�ů����3�"�H<o��i�8^m�,�+�g�=*#8Vs�.�M��]�%�95ґ��;�yig�1�
���}#\�|{87+��'������S3���/�)Q��n֫�T/����)F��[�%/�8L��lY����O��x�N�t�v��k�jzM��4���9�j���Š��I�tΟIevm {��%4�"hU* �}���ƙ'J3?ÿ��f�n
Nҡ��]j.�`���_4e�?�GLlk��P��\��\�<\������Ckc4UU�,�\�v�$��w���X�s��S�r�1�Z����p:�=(��ͺ�T2"׊v��hq�K��1����F�k�j��E5���t
�Z�q�}�{��"�o�V��$�̜�;[�s���s���󙄔ส[�G�����H����,��4h/X�z(����4��K�q�3��5EhY�9��&m�Z�#/M����'����UyV0�x�p�N�������یp�:��:b?����X6��\��p��_U�|?:FUd:�Xh����G��N +�;��AY�r�?���=0��M��q�}�V#�s���B:8�����"-���OͶ��r����!���:!�'&�bg).��B{��!���t�NPJ�[/�"O�p���a���+C�̥>v8�х��cs:i�C�>=3�z��t��\QU~��#�.�	��+��Rk�eΰN����4	_�!w��$���EǭP�"��sIw	V�����}��L&�l�޵B,�X�8`����(�ý�vl6�]s*��g8�?�u/*J����d5Dq�[�t�05���H,��J�:{M/:@	����3A�+�l�c�SێP�XA&�4x��q��'�Ѝ�D���+&gB��i�����n���b���c�U!�#�?��9��a����l�v�5ϜW`#�J���H�Oo6n�V�����)�wwI��c�*��������+_��Ch���t�l���%��DC�"6Y�A��$!�$��s�6���O3P�����{�?�$�Ő]����SH�q���~���H������fr�JQV���1��7F9ڤ��+�����"b"߂{���2~�&�g�䃬�Aq6B��7(h觼����:ПA?���aa�OhZ�IV�TO@X3�[ŭ8:zQ'�����K�%���q:��X"��� ���_�C���I��U����:?H�"�xiso�l���O�0�j�e5�Weδ=�,���z��orh����#AK��p�0_�-�o1����xM�Z�ö�����\YԬU�R���;u^�L'|���7cݏ��v��TF�D���'�f��ǻ���`����|U,�w�����ڬ1�J��.�z�/ hP,�5}���8�$�����|�m���q�c�������E�y�9l��5�x�=�)ß;��?$
 Gv����-�ژ�?���Z���
6O��^��o��睼p��������]Zi���4k�ӁT;�`es���&-���t-��y�*J����
��A�>�L�.�~��!�	1_�5ZB��;b'�
����[ˍw�B�3��(�<6jG�t��Ե��5~��K��{Z�T��l����S:��o$yxo Ʊ�7���Ja�c)ܨ#ߤjC�7m�>y+�Hi��
 S@[q��Uwx�^�`�}~����D�,�!W�j��f�L�z���&�h�`���q�}�����*�3�}�sE�vVU7q1��|j�wo���P�v���[�g���5�$R̘K
�����a�5�6f�����^W/����t j)��e�9'a�8�~��׳�P�6���}DgW��V63K�3� K�=�����a���V�������R���A{�)S�������)<���+u��1��Ą:�|k��"�����'��J3=f1���w�2�fǸ�qkV6�m�j��� �-m��!�����5����T`~T^���&��{��
��@p+�����vw��j 1=�Yb�1�\�lC*�;_g�}�
�qG�ݠ��^��$A5���"VRWX���,�0qj,��޳[���\� L��J!^��	��E&M&��C�9a�Ƿag�S�1�,K�q
�1��r���yuZ�g<O�	Y���hc��W��n��*����J�bSX����|g�C�z�������0���� �ۤ����V1���A��t�ږ࡬	�e��#z}��R:S���Ε��g�E�ɔ�tY���ƏP[ ��m��������ɟA"��'×"����j� �O:h�xc9�>�S�� �(a�I�w��U<��G�x��7�㜓P�d5�ߏ���s�M���w;��ٳ}p6���(3�\$�́���e���$�|��] �
]b'M�x`�` V�-���0^K�"[��9�8�`t	����W�����ٝ�$h'�*d�5R�Z�ý�M}K��Z����~>YܠF��DEWo��Q4U�d��c���b�^7�ձ?*���	pG��4�M���Y��U� ��8 �^r�0t��HB�����߰�{v�m�r�8�Q�:�T���z#H�Z���u2\�S	�}ts0�O�`m�_���DJs�~�nzW�Oy��߯ߎ�0�:X;��{�k�?\�NY23��;����5V̍`�T���������2Q�W^V�Ci�C6|���L�49�����l��O�����f,S�qO���Y���dùlU���[�S)��=�m�FZ���|����E���`�'��q̡��~���nK���4��3�3d�N�lP��9'���eW��4!f%�@9�N}Z�ѯ�c���6��,QTΡ⡎�Y�}���:�l!'~��$53&W���-�E��`c:Z^��3�M�'Gß���x�97�#JV��z�R֏���'�/(�$L5���߰6�ˏMw0���C�A�KM�q��Lo6��,�{X ��Eo}(Q���Dd����S��u�UA�F`�NBs�F�N�8[qb!9�K�^���(�h4�;�Ϻ�6���G{L	�dj����"�b�5v��Ԣ0�5@���2��^�`{�c{��V�n��V���ڴz�F��E&T�(Tap95�������c�U���):0�{G!�i���7>dJ\��=`��چ��� �L�ۏ�����W�>oa�[^�7t��?�Rѥ���+��0馍,���!���d ��9LY�����"Uo��q%�	%���}r$�|0G{��l����d���Z#������oX�FM�m�Y"���j�R�<������}>�DV�L*A�d�q�J���$D��q01C���]>tz�E��'��S��p�Hׂ�qe�h�@v)L��L܁�_y�PC%�YzK�|�G�V�j;�1-��X����aC͓�D2j�~Zoe#��be�͌�3O��+<����2�>����+ʗ�s��}�<���c�&GN#L��{j�c�3�<�4�U�A�0�0r퉏�����E�£S����d��714��D��U���R�@&tC·�;�u�y�	#�}GA�=�ϟ�����V�a�4g}gF�m�4����|#�U�JY�!/D�(լ\h��żBHY�jd��]��ujD?�E�qv,��ҕ�[��
x(Uf�ю��H�
��Az�8�����iI/�:�/}at��*��3�bP�q���?����競���������8�nx՝�#����(.� ���=W�U����C��f �
<�@�u@���H%r�� R��r)V�1��
������W1����0����������5�A������{dQ��s� � s�R���lF����BkY���*˸���U���H�܋���C�K�~���h e�4�iF�����F
@VjWl�����ꃩ>��}���]����bxΪ�� �g�%8�آ�U�`�<�����!~��l�׶��.{#�=F���M�Tf$/1u���I��'Aś/PC|Q�`A,e���$�#�m��=����K�)���-���i��F����"����{D���|�%W�Y��k�S�V'��.U��pq=P W�wOoU��-u��U�x
���'����w�!G�Q�!�w�����9�K���Q3o6ԝ�q"�(�&[�r#lAP���L\��Y�}jjEy��QP��)@�#���F���IW�v����x.��ל��'��ȏ8T��j�d�t��Nr��_��su�%T0��զ�<��xFy�뵰�^6�~�ڶ�F��8 .��J"��8h�½�p�E���Y�͍>�γ�j5��)�0>�x����T� ���p+��Ԟ�5�Sre&��h�b���N�u�[�K^��t��L�ʹ��Fe�:͊��k�@����z��ۂ�̩��}��+�N]|oxhk�Ѓ�F�.���t�D�*/��t^�Ht�p��S)y���n�1g�	q�o�B���I'P��b�|}�"5� �*=]���^(/NCC��ʼ�!t�0�K�=���/6	q+�^B�R�٘�����B1�gF>���T���C`
�y�(
���B�l6X�L��y��a�5Z��n���#V	R�kk#\�$�`B�T=�^��Fz�Z/�[k:�\�����0��qi����$ɡ%Vu�OC��jzj+�s�!1	v��=̧�Б?���Pn�C���G�\=sl{y����	��B��X~��K��Riy��Aple�r����;�E����rjVĝm
��VW���ҋYk{U{tָ��}I�0k]�X��!�Ƀ�1z�^r�
��T�3���_ggg^2���4#��,ln��A�y>����䣆��Y_�d�ϕ��h��.�	���JyNa��'*��� ���#jk�L�����P.��4��&��橤����!@@��46g�
+�����SN��#�f��W��ɯ�����d���n�F?Ì>��h���=lE@(�T�2��F�D¶It��G���RD��p��.�2#:�m<��,�Ď�hd���Z��is.��Ўa�iLQ&`�T�5�K+@��W���ta3"pME`�vЙ��jʁ��8�B?(�hC׋��w��hr� Gؗ�E=T���i�������aȐ)�5��{��6gw�S]"a��?�K�2)���.�9u��efXih\�����*)�x7-��;0"R����N�+�l�te���	��7L��:����X��gG)Kh��|lY����:
y�%J=$h~���&�)��K�ݚ�g�	��{�����V[ķZ������g�;��~�C�O�C����-���8��43B享]������Or�u��qSͧ�'��Ѿ���W&�Xn�gP:�ʂ�$d����5�.���6�Hb5���ŝ(t Y��95
�w��Ӂ�m��>r��U��m�!`,y����æ�m�9�����k����ډ�!��%�DC|]�Y��CFu���sE2V�ӷ���%�R�ImU�`�+�oi�T�QP=�/�V�|�dT����B8� ��"��`i �ষ̕{�xƑt
7/|.�0ܲ���󌟶��)ܰ��&�\���P�$�� �Uo&�na'��_��/�KÓ�i��uO�cX�]A�֗����]s� ZH��?��S�sd��p���ɯ�ǰݚ�t	w���H��J��H<ָ�A��R�^�$˘e��#��A�i�;��� �>��(��\	��_w��J�HH�f��rʆ �,�N��DV���[�QҚ�ĵ
v�5��<7_��LW�"��́�G�&r�i�k���( _cQ��d���rh#��K::�l�1���/lw�.�̌+��@@]T-�� a�~j_��L{�X0��(f��1�(A��>A�*�0��	
�J��J�g��+��߹��t�:,�a�W��%J��4���MΥ@���FW�awc�3͟A�<1���;]�
��6�0��Z�_~��VX���֙ՄK���:sϒ� X��@8�  �O ����5�s2":ѧ��1gT'_���M����p��c����E�EOL���*��9p�+b�O����N�@dFR�����
~M, OG�ưQ J���/U!��N�����P���08�1��-���s�����+bQe'L �g��D�ZGAN�G���w�>ؐ����I�o-/�����]Bf8�����G���
�@��z|�f����R�U� >��[Hף�MM���پUg�qi�}G�ƔKBm���{okx���W�m
��})� ���8�iX��z�P����_T5�_[��08�ù=��fw�YWs����������n��.�b�4���������j#L����c�VQ�C��t��.t�h�[�'Q�*Q6��EwA���T|�ɩ ���;�P6��;�݈�<ò�+ږ�PE�� �L�2v�V��ۮ�=~�R*]0��6���N�񄒬���I�Lu$��]�u�]�dd�����I�v2��C4�2G|��zI��I�ȒP}`)�G�lf�$�]�P�q��=��K� �jCU_���r9�U�(ȿ�hWa���¬u&^F��[U�XQp`'o��+(����-�݂�QT<=�`Re}�E�g@���{�?P)Ѷ����Yd|���g��'���C�OJ���q���>���(��0.&,���)28�sX?����ެ��Yf�����`�h
�����y��� ��?39���R+�`Q��,���U��O?i�@�E�Ёo�j������B���M{�;�Zm�@ca�d�+o���B���[��!�t}��i;=�\T��0w;౿`��0��ƚ< Ub-�eQ͒B$i����n�o0��2�&��WK�����f�Z��̓2���Wjk�pKC�#�>�K�m��A��š������!p[L5O1gry���o��1g��MKwΥ�Ҷ�.���T�W�/t��<5�(MtHўboo.-Y���P\ݧ�F��
��t�v���Ѯx�.�
�~0�rt��wc�����6��'����=3�~�ٴ�m���\�0| $t�z%�M|Nr����cK>d�l,�0�����-�s�����<�PXa�M��S=W>��Ц�Y��@��B1Q�#�ʞ�Ҋ�.���V#�"Z���B
QF_*us��1Z�9C"FZ�"��z8�-�'�X��
gAt�js|yZ�Kh�@sٹ�uxh��p�=�=����@��S�j�ͨ�y4\��A���A�X��Rw�WwDC�m���C��Xk�sJN������#l��uǦ���gH~�Y	xw���·�{�@��ɥt8��ׄ[G��/.1�#*��W�\����	�2�WJB�o�YnP:��3�L⥹�3��C���Ҳ^H���)}�A�+0EL��\�) ٻ%�nB�B��T������2Dt��n)4����w���f8 ��ьֺ����N,��~�.MhI���&��͠YF\{V�m�lو�ՠR�>����+t�ˊ̛JÕx�r��҄fP�`2 ;�en����@���[oY��Q8:�q��e��+�;����t+݄E��m�c]z�I �FƉ�SI���"	uvVq��4��������>;��+5E�K�W��F���AlW�4�9�:$9b��W;�03^�̃�l�>};�S���A�E��|�������>ʟE��i�֔O&��O{����=��8m��9R�CK/Y�'k\�R��"��in��M	��=�X.�6�r���A��P�����ͥ�@���>�o����W.���~���3�-�(�w��J��C�%r�ܚ�,%�NOd�84a�������\9㝤�6@�2�E{l	\�\�%ʄv���fYάx�*>�H��|�PR?��iG w���s��8$���n���a���7#��1��5�V�>/⤆MKa�v���Dqz ��b6;�������E����zL����+=�^Uo[�����7�()���S��&.K������-�kt`���.�~ذcҍ{��K7�<�}�!̣y�0��sejK���Bo�p�{DR��6l�ܻZ�����fL����R�W_A�����t��PF-N���j�T��RY:����\v�����x|��*�����D���(p�6�BZӐ{�n��)ɰ���PwMO�>�> �E� � ��jk�J�Z�4]G.Gn���题a��դpFjj�R�*a���Z3dY�Y�%����܀ebۓ"�`_����l/c�<z䣨Ȇ���(p�e�(���Z���/�����ZA=�9?���������
���ٯ��ߓ�X�G]`\�Ӡ`yD�f�l-a���T�%x�W�@h�_^��nxT7�j4��\�>E��Wn��q_Y���g�0\�Rkl�x:%��1IE�dG���^d�����8��>��H>�-�=��}�s^.2��	k�&��7�W��ǹ�̈{�b���
,�d��U�c�5|�kR��@pX��cȂnN�0��L7WV�i��;��k�}Y{.:5 ��d%%R�
�)�~Iս`'3�wК���:�T}[�q�=w���?�
�)#彠������N�A��]�.]L���%��qz�x�1��gH��xĐ�h�4Iu��O�+�:>W�.�o﹒B��R5�� 6XŨu�j��WзN5���P 6r��%�97W�Gm�&O�{rn�����F��0�0�@��=�GN:*�\���M��ŷ�� ^�c�m'�r�
�bۙu�Z�*��C�"�9iv+k`������������|o���7��=
�@��:�~�ɩ�ͧzȆ-�n"ʝ��&R^0���� �g�5����[ϼ��3),Sr�$Xr0N�u����R���3�h�%@Ǳ�7�r��K�t&�~�rL|�愜��4�ѲE=�Ѣ��2�pΫJJVX��*
���� x��^��^�p�%=���\���A�aQRڝ��~���H�LK� "01��pu��fO҂�]�-����ڗu:ָ��X;t�ժ�<��z<f )͌+[ט@x1,A�]tK�%$������{jD�5��_Yps���F_�u�;��ÁEV��Ĳ��X_��@��hˀ�f�s܁��~�
Հ�]<�h��صأ�ژD�j�9Ҝ>�L�G�qT�����M7zj��q��|8�n�Ꮇ&HIy�kL(C����:�^���|)�7� ]�J|ح��$����s���'�{['��RU���3h�z2�����YPV��l��)��Y*�յ�i\DG��L	ʼ&&2$��[�Aa�g2w����Ċ����U��ERer�XB�q�0R��=�[j�����S^��=he��/	���]Ax�<ąI���~��Ŧ�b3f��#� ��<i��vU4;G�Vם�ˀ�{6�(b�^�Y͵)}lk�Dp�,s��Oa3����3�{��H�L؏����P>Fi�3 `݁)	�pc�"+�F���O��rdV0�ڸ���
�a ��G�݀]�@�f�a�l����	`���!����R�d)�ʹ�0L��:+`YX��̈́
�� �DQϚ&̿Kʗ�8���g��L���~��:`�QMBs: ���;!��r�9�)����Ao�	�:�Y�v��؝��p�Q��!(&g�!8zV���}<��"��ak��X�&�3b�p���M��;Ƹ��Թ0%�۞���,��Q���f9tv���c����<���y!;�:]��2��o��W���O;�j2��E��$�{��WK@�o[�H^M3�C�Ȏ��|rv[,o�N2kb��{̊�]����.�G�C��	-݆�	y��K�_�Fl�SV��j"���U.���IM/�y���v��6/H~�'�)EBb
�uS��K��U�Uc�b�mHŢK��ʡ�6y�`��<5���o����P$�l��vL�-��}DN�Û�:��#AJ�R������U�G1��WK�F��KG��2��u|EWL��'�IP��m`���q��W�7�,"��r0I��z�V\��fJ�>6�N^#��L����#��{�M）��3�E�;���3������F4<W��ʸ�W��櫄j&3b�+��_�X����V�=v��kQ6
���хt�Z]��`H��v���F	07#y#,?�F�W�Q.k��~i+�|�X��탧E.����FZ�ہ�p}�Nn�XkΡE
�ہoG���`�.����I]�(*�6�sGeoe�[��Դg�ڀN�5q
�NN9#�ЦO��Y�A�z����ԋ�X�{>2�ZC�X���^�ߓ�z�c�am��iɢ�xk�Md��
�5XoO��׻�C#6D�6�L���Ȇ^0=�P��=%�ÓCy,V�̬iN�_5���N��[F���x	��G,��޶�^�uh��'�ۦ���F��A�Ã�"T�&\[��������% m�?���y/(z4�(����} :�{ �6�{�\��,�舘�y�J��?s�ϸ��&��S�#�2h��5��c�j�1�ޢՄ��m�1�)��XO�8Y]�J��I��z���Y�Ng�{
W%ApN�̀p�ӖP���'��\���K�sOuHO�HWԫ��W�)x�W�2t{�?�-��Q�K�[8�r��`�����P0�=�{�lLI�f�ʠ��j� ���0��)Q��n��	g7|7�1���}�W������?��,x�,6%6��+�|�6�ƪ����	՞��Il��p���'|�Ǖ�B�<��vD�j���SwI��B�q�2�'-�R+"L<u������P�u7;ĝ�z���'����J�[d�sdc�eK�k,�ٳ}���[�,ʇ�s���a��Gu�g$��6�ٴ��0OѰ�v
��-���VM����jz�B'�&8I�cd��_����]�~�Hͧ������ᴨ�8)$���L�V4��B;�<���I�J�*|���Y;
z��<9��E�Gw!�c2�كt��*���g���*��7�S���qn���ă���:�~&��{%���X�)���v�2��-KM�P�i�S|�'~
���P��46ak���xr�pƣ
!K<�M�ƕZ��j���1�E8�1I�U��ZL�ȡ�RD
��~}|�hd�ݕ{gc����x�A��g��+R`��s��0�65��c��|��z��s���O_����
F���7he@@Y�8[�Q��^d���T�%Y�s۫:׫��R��?V��b}33�l��cqr�-��H���`�R��R	�nJ�/o��%O6�s4�~4�x/X�4�V������ta�BWn��X�s�R'U�R�H�8
H�Z�S8Irv����)#h��8��W1i�G�5P�.���$k0�s��V��G��o g8l�JB:ItG�=��lL^�]؟�¿)��C�
�t6���g�D톢�O��������48>?1��@�Z̫�z������d
��p�q�F����J�z{���d�}�M	}�k��a@����Y��@���7�X�{˝x���rh����Fu��0r�}0����YR��o�Pc����e�;n�<���ݍw�Ǳ��.���@oUt�K�����c�x9����C��P��i3]��9����h���)��͙�}.��~&�P�/H.9	]N�2N��y���?�y�"����YOT>͌#b��3ŉ�=U�x���x��"��ڻ��upF���C����\�6֎�۸����[�n����0��!����R_�,&b���6C�=i�����,��\�Q^��� 7�ea�@���]�$��nȮ¸�4795�<��"�V� 0>�/��6����sŸ��-�w؋��� Qx��ӆC�XW4�I����)J*��Bzb����Ym{�^Y�u�Y�>���4 I���n˪?6W��۱��f~7EQ���4E_���W�i
�C9а�կB���.t8Qx��ELoM&�a�i3k� �D���N���^��=�-������Ƕ?~-&���ëxi!)Ǧ���&� ���WRַ��C-a{~��ۮ$`h'��?�k9~��2�5ԃ��kY���s�'&g�Xw2�YX_�����w���É�
�WQ�=ٺ|��3�t�^��QMwtC�2�+g�%�e�A�*��9���n9y�
�G���D�+��*;��NTG�`2P���<�%��6��yh��!��SB'��������&�v����K�h�.��k��;��a�=�ѽ8F�Y���ܩ�T�@^�����O)[q�wn;B���)���ڔ���9��l����d�b��9#E��I��<{�R���[&�D���N"�B�(_-<�x��.�a�\����)/���n�
ԄZ�!��"�,�C�oq����ю�'�6�bei�N*w��Dp9Ik^$,�|�K$�����Oj�}
�!҉�.�9|� RZ��Q#4���g�Y���j5��ꗫpP����|ƕo�%�M���mnԘ"28ϐV��#��5��N���ʙ�Q~���ͮ����%�.oӛ�^���N�Ǥ�;�h4�J^��Cmޖp.+��Z���s[���5g���>ƺ�u�1�J@/W!6)څ�N��ߟu�����N�C�jvu�B��EL��BĪ䨤�Ur�g�aL�ԝub)^���ш�O�'9.)}�VJ1�nO>=yHB���Ꜹh@����E-���2�C���3"��(^K	�̙1�>�Z��ޑ�(g��k-��W�p�YB�ЖA��s������o�¦M?��[����I��$`�o�JP�9�}���#�d	�N�Ԧ5�l�@?�c[��jY�s�oG(fLs���γI �@�L�����V3�i�U(+�����?�r����$���̹��
x�c�A����#�(���x`8�{�pR,�I*GI�󜩀��+��\v[A�+V2e��ZC�S�v��&�!}�k���d$�{������r�K���u�;����O������[t�]���uy	�O(P2=]WN熿�C�B�V���c��H�͆A��/l��� �?������}����V`�½o7�g�[�(bю��`������RK`г#t�����Q+/���A�|�4�o��u�QTKuh)nl��	i	p�y�{��.�Q����K� ��ܼ���E���`�^�eߔ���[.B�+��e���8�Qt��O���&W�L�����8!j*i����v^f)�e�l�Ԉ[�}{>��R�1<:�N��+U����7�jk:$7:4���á�����T����L�q����sV�E�i宊�;�E$��6�`�4��|`�Y&��=�r��!o�4�q�S��AE�<h6��&�������.	�J�7��5[�JQ��IE��"�~jw���+�����I������;��_�+LPp`ڭ�7�=�D�Z�ו?j���0m�%:]H��*�X��)DyW����L�|����kE�:|^�?�r������|��!�z�D��%3��W�Vt�9��G!������K>)��?O�Y�pH>:|`�ub"S�y�(�,����R�ա{5ݿ��sXrsS$�ųc��'�4)}��0*�P�Mo����>�-�	�#M[��0x�z����*���a��ߥ\vr���T~�ѳ��}�x��0:O�S���t!���j��y�wĩ"K�d{�l�}�c�ʹڇc(l9+HE6f��fa��3:�ުN� �������fZ��8��(��IQ�w�ۥ����O:-[�' ��B��zz,�r��,v�r�d�3�q���b.�W�У������{���Z��)�����ן��-ط��m�M����ʃD��ZI�M�O�p��N]���º;��+��Y�^�W7��NΓ��'�ӥ뛯��s�v�ja��\�$K�00�%*Z���鸸+DDl�^xy�O���u#ĉ9��HҎ�����(�I'��ݖ'eV])�۱�?W��L���<	�*m�B�b����k��~}��H�F)ת4�c�*.4��@�gl�a
*��MT��Ƀ�G�z.�����(b9�p���;��/���ɢ*[oI��Z|�;W�����gN�HJ���r��p�?�
_�e��i)ңi��Q4��&6��r�C�
e�0��E[���
|�F��^�Tʬ�怅�@�����,�kD���a���[~�oX�Z�tT%�!3���̦��Z�0��.�K8K�M�	}�o�By�o�hF�� ՜�Ώ�8mpS���S�֬�)�b��V��Y��?���M�f�g-�4|�����>�;�м�s��.VRwO2��<��f�Sq.�pS��A;.���L�R<��W���&�Ya%k:�6t��:o��}�v��Y��HHƨ�4��T�8��{@����R��!8\Mf��
0��-��Oe��PK�$�]�p��<�Y�L|K'[�y��0, e�&\�%����	��࿎_�-G�����s7�������.K���iT�ᣙ�fvF0�O�)�H�\Ӟ��X�޴n Zi?ٯdE0C�����-���g�:8�j�{4�o���%G���um�Y,~����SΙ]ř��]�>r��β��H�G�7�6��ƪ:�&�ߣ��@TeK�a}�13�ni����"��XOq`���e9��ln���h�GG� ��E�զN�~�1nX�_����(��%e�J,Ƭ樍���/���fԽpy�NY/�9�m�D��g=�� p�+d�,����o�ւۍ7���%�9c��4o��a�x�>���u$�3F�@Q�U&+. gQ�n]lYeo
s�m�.`1	�?��d��'Y�^C#="�O�I���#+=�R���%�E�_���K96dn�?��C%�
�9�Y	��$�$���	U+��!���'��z���\���LE�4,inV�t�t9�~���������U�G���kJ��!o�O�̭# ��Bl�����G����2�[@K��p���J>sτ�OP�QF�+%�b�s�vXG�'��;����B�U�B� %v�|�W$�<@KW�E�fh���p�F�!�eO�����{8�j�yH���`$&��D1��_��}���t!*D�t�=���%�j�����6���w���&�{��J��M��� -�'_N���.<��F���R(���S�����< NQ�;>��)[�5�����;H��)g�⥼�E�̖�͓>e���>�ҷ��J���X���c[��uL�&_Џ��Ȁ�R8nh#N&=�/�f��Hs ��Sމ۫�=�Q����(��L��*���H�2�]�׺�y��7xIW2
��C/[�]wKf�<;�m�*eJTB��2�3�gb��s$A�T��0�o��	�*eI�y �(챲ce�Z�TL��9���@��'8��w���Pt9=}����Oض�����x���W��c�V!��k|��֌'+T�c|�#�����n =�^�.��O�1pv�4s
.�o��[ò+3�8XC�{���Co��4����L�x.��/��kkp��*#�c����E�������º���F[��u. J���NK�ᇵ~�=�0�lou�$_`g��@���z/�~���7D�-���J�e����t<�*�'s#2IS� ��jO]՜  ��d���u�`�jg	�Ɵ �,�X44�3h���ے+Pq"(D`��XJ�+���:���b jW��?2�v ��fs+��9I ok�>�K75��.��q�U=fT��0���ib�1�� $��/.�>�%'�*�:~��c?��HOJ���~	��7�p���g��F��U�''�8�1��\m�� P{a���D�m����p�����f�߸Z�V���P�ߔZ���'ܒ�!�1;*�+��J�?3k��Fᦗ���dS���	�7�nH�D�3~�ܼ�6Q��������9	A�>�Oc����۶��/غ�T�摵vn63S��At��1��Go}��}�2�#j�ÕF"�^���8���������ף��]��wK��h+/��6��y�c� �@y�q9�� S���̞���t����}1pҞ	��+�,��;f���kxzgc_�'�uvFI�-���Ҍǲ��-��A�u�0�zĖl:mBY0�����Z����wQG�o"�:�WN�f�R��I�s̍h#����I˂LM~s�ke���Z�����l9�j�٠0Z�]���ZK��\�"�@#���Kڿ$y��3���'"��nG~r�nb��9_���a�Ҿ��������J��:Vy�K�dx�qں�������R�z�`�)�+���Ӎ���p����®e�s�1�~�x�����j�y�p?��j+�G�3��D�rdO	D�;V�$\0,����y��"NJi��j��zi٫�̭ܻT��--���k0q09�N6�s�<G�P�.|�pf��ם��2��d��҄�O�̓$��	�fy���r��(	��sN�Mc��Vܰ}"�7�ǶW��/|��| /�c���}�muz��TsL.�,P��3.���Ga�{����cL6� B��)��J�����	��0�<��6���M��n�b�N����O�b?��O
P���m<ю�)��� � !�өrd�o����7�y�x�kK�����d���'z�~���eh���Pv[{��$f���~�����)y�ʣ��'g�:Bb��4�^u_��M]�:��_� 0��ʹ_�H�;��^���\��C6�����.�n�NTO���ݧ|�	2�'<s�[��	�\��P���N��l�B���0���򩮃�'�8�"岼���ߕŨ=Tn��X勼r��R{{��l�7��Q�o����a94��{hol�G0���g�2kV ޞ�kj��Q�͎f����5C�ߥm'2 MDG���H����mf�⎊kjҚČ��l�pH_i�8́oČd�W�r��(X3ɊrJ�@]��6�)�Ͻ�_5xڪ%C`�ٲt�(��o�����Uz��U3�������E���k�:PēR��Z���<��F�y�����ˢum�z�J��Σz�����[���'�-���
���s�5�{j�E��6U�-�HN-��f������C�;���/_��p���S��ۇU�J���nq�2�������x����Q¨$�?�6�Ai�(^o���7Y��	�W޲��wL8��KL>v���^#
8�&����oFi�T������r���9?8x0X�d�tiv9Χ��cH�b/G:�S/�#Qy-K�Ű���=M�InjjNv�ELm�s��'+ �0���diw��O�{T��������o̵Gx §��]��n1��m��G7���"j�q~+Sa��+�?��U*�Y���Sv���f@��֣x:��<�P�3d����������d���dG	�V�Am5]b-�bQ��T����u&'���v�V��M"C����/���nޞ�Z����h
GR��[�.��
}/�~H6QD붎��޲�"7���� n�~=��nE���T�@|���M+���U�����tn���ߋf%�kpk��O%�VU�RH��D��y���*U�gـ[x�� @�R!�2o�2��m�ڋ	�q��3���=���T���r�s.�\�^�1ո$��NO�$+�� ��XGU�{������C$��]�
�:����C�6��u����}z3��[�/�c���T@����||:z!� ސ�Yhh'�(ԏ��;tx�G��4��@I!�l�Z.�A�;��hL;��"ɳy L�H�3�N^z�30�l�v��͎?4�p
p��ox�����t�b� �����K�/-�S���@�	kX	���傔m��f?6ZA��C)__g$�]:B�y�t>4�Y���؂S*SC�'@��󱧪��Ea�H�׳��n����45���3��]�2�/K�G)���dzǵ��H�עP���VM%�~�g���'���(�t���҉�<�V��0�?�}X榩	��{ngR��Ck�ȟ �ok)p��J��f�j�ͥ%���:&e_`���?�@.6.��+���+�&��UX֌��XQR�fѧ���ƛ������u�QW H,,F$R�6��{v�'�/a��j-p�x��&#v�\hf&��H�&��1j���3�E��jq� eI����+-t������m �!��B�*�]ǫ��=��
Z N"�Xk�H��xA^ߓ��>�>?�V�����b����UD̽:�$���������n�EOi�B��JA���ڲ�C�|���/^��r�g�X��<��آ�R��
�<R��>|>w|�, R(R��"�M�4.��t�b�e��;5K���-H{W����~�/@�om��!�s��=�`2�e���@)�W�{%���o��y��tLM͢=�`�'@��$a"ŧ��YD{I:�21��$�A�#C��1Mj�I�2���%�\��*ꀷVz��JE��O��?��(�{���/��g��H]_a<4�'ı�^&���0�E��5��.�O�6u$���D�n��-@�/Iy����Tj�796G��H��[|�&�`�<)�3uwe�����4��:=cl۔�{Q�>�i�3f��ֺ�\b]�B���Q��z��D��4�xY���d������Mܑi0Mt���5�ޓ�������V�~����3*������=���%�d�#������%�X7G�V��>Lź4pAW�IovR���m���Dz�z�N\�v��\$l���(�l��v�P	��%g�F C�G�';���?�W��(v�k�N��e�41���oL�e-�U�&����hM��fӝk��'g�C��{.��.4������$2O��6��FפzH�q�
>.�㍰&���g�Sѵ��w������7���Q��+����Å��)��t�����" (�9����v��z��=�	G^�R��R �P/%����l��[�����[^��ނ�˸QA�,鹱^�'�S��dӀ%b�=�=��e"1�pr"йI~S���ąv��?�z�R�<_X9��"5��*fjD��F<�ctx�[�4�c�~�:�_��NN�u��FL��qp� ��[I�I��ȷ��%L̽�\��B�TLQ�$s�派O��!�ӆ��,�wBx\�Q��W�_F.�+{I���*pc���h:h��5������T��sJ��@�s&b��Z������v�x����v]DT����_I��<N"��L�E�Ds=���n��B�:j�S���Z=�6g�%v.��j�>^�h���(�BDJoF6�蜞c�}OWr��w�4�\��Iݙ��eO��WC�qc�Ñf���(�:�|_������!�7�
�_\e>J1Z��y9\��8wo�"�6؄$L<��5�9I(>@�-/3y#��*�����b��o�-����E3K��F�湟Q.�CDg[�r�<�������'O�-���	�i�$ll�n��d�G�Sv9'���������0z�$$Æ?5�P�X�Ρ��(�i��_1"�J:Á�n���}ŌZ�[��
'���fL�OLϬ.d�x��꣟otyR�ƶ�3�[�n3@����'�N%�ǳ�R�5��-gV�����+t!�4t�ǓL�a��=�H��k�bF�Gdɞ�nH�r��*ǲ��.�k�I�C�b�EqG���NŞ�����y%Tw��~�)}�`���l|U`t8 ,���^��!�~^��+Մ�JV�"����2jU��|��9�و^���(���8�p��㗬O�c��G��=d�ƶ�F�{yL��Ǘe��sەHԂa&�����Ȗ ��5�7�v�pнāt�6�?e��Gy��·�Z��$[��}k�%����V7����g�B�Op���%cJB%���%�z����qvn��$���t�2�-c[���4\�v��'���㬯XY`����u�(�E;�'a�V��Xl����JJ�0N�Z��q'g���:���,_J��������α�����M�'r(�;"��)���TI��*`w�qqHy'0���*�E}
�9�xU��2bd��cR"<3�*�F22��z�|)�5��E�\��_��&U�r�����_�t���	�Iz.���1���],x���K���ɺ|7,���A_{������9�۟�v�ە���;�+Qfq��p�rړ}/WV�[�F�ͩIK�������M��nfL�S������%He�%�}�r\��ݒq��J׿���3���^A�'�E�^���J�e����x�o���\;�{·���S�����4<�Z<[>OG�����g�.����
�	a�?�@ު)�����la��S���O�<�J_�ĸ�({8)!����EF�u�+�l�{�d椗����7ca������Xj������"@$1�d�!����܄K�NqC�=
�/݀ߒ�YÒr���ׄ��,�r�.>������Ux�-����)�҃�f�~��A�I
l�yv36��%���<��pFY}����?ta�J�B��U��3D$��*:c�7Wܹzc
���O��� ����7D��/6�q��t�og�� N ��
p//�S�m�SAʓd�TB_�A'���|�5�W�B�3ڿ"��4��E2��\SO�'�b�)� �]�`Gy�c�;az�9?�xr�e�M�1�
G���-s�ʓ����=���2�o����{e����k�jz^;c
���}Hag�9��g���ڍ=>�)�B������~>�g��%}�Z���Ni*�x���ѩ(�+�|W៝R�FB��i*^��>��q�	j�{�E�K�J��¬�4�]$��l�L0kή���� ?t��eBVl�s6M���#�?�ٝ#���)�󲬇I�~�:���U	!Մu�N� �U���W^U�_s��Ћ��W;c'����?$�e;�mK�+���.�Y��=L�ړ�̶v�7xM[Ͻ���"�������q������7oi��DF��ƞ�U,�uX�W��DV�^K�V�'ϋ����ʻ�}4ƋT�Ѣ9����Qv�r'Ń�^s��!*(�EO	�k%þL�a&���7�����0 �������i�Ǭ�;R�E�V�b.�8�MH	�����S#����jWW�u��N"������I/�d�����t�Mgv�-Y,66�������wD��k4~B$=Ĥ|�㑧 �*1��1�"ޞTe�Ι��ة7��]����Pk#��J�w�V�	�a�z��� :��c�N�Md0$�<�g�����R�ݲ���W�e$3��>��0�^B�G�ǔM�����ǩb�%�ד�H�����d�[r
�Wc( �
(}�~j��#����m]#��ֆ�J���G�N��^��,����T�8�i'�b���V���&��:��������9d>YDgJv��[��*���0g����S�Gc������@ִ�8���z��.$&�������k����੣W���1#¦���o�$^���9'�9�oe�yi�HZ÷ʉ��C��)g��H�z�ܪ;9}�� w���֫�v
Ow�xLd�c�x��!V���Dh�"Mr'�F4;T�]u�F��ڒ���"��<O��X�RL�}mS�|����
���Aϔ;:J�Gs�{��HɅ���O�q6|Hŋ���[�W0V� �������y������0���=q�����d�	[[�`!����?��ƪy�:jsB/��1{W��t+y1���C��?�Q:�6��X*��b�����c��sn��h�c9]���s�	��MT@�R��/ؘ5�{�#���g�֣4�y����r�o��	uWّߜ��?�Ƀe>>k:Hz?�H�0cӼ�̵s��+�W4��h���C���q�d������-fDYeN#AN`	���=|z|��Ax�3$�c���K���(���6�+b�*�y��+�	�_�MMl#�! 4��^��C+�.F
���B뜸���"_M{؃)��iz4��=�_N��dF�F2�>�
EYh�
.��8`�s{��G�s��j�3:Uq�j���#l�^W���M]tc��� *�{~I�o[�ݒ�3��g¯���vJAH��S��R+��@�c��ZjÞ�	I���e�'ˮy�j�>Yӯ�w�U�jG�<�V�^%��`l��F�����n��V񯵛r�:�%���6�'���e�`#c�qq���_��T?37�Nʖ{p8"=��N�nk����@�{�w7�h]g�os�,�T���l�ʤ��1Uo�,�Wec�����s�o}"�S!2�S�1���!�����8���߈.[���e{U����P7#H����}#ut��Vw�Y~)����"�I��4d�>q��v?
y��D�.[T�[���e,8�N9��k>8��1��D�������9QU�u}�2�}X��M/�כ���Ytܔ�>��k3&��},f٨0�!�E�`�\&�K:^���鋳IV��9�t�K�By{��0�!�#!�6�W+w��}C@�F�֧������8�!�
7�Ӡ��ԡy_����K'�#˪U���w��m �*"��HT�Ӳ)�<`d��dr���Q�!Vra��{���ϑ��{��J��1E}�3m�x�;�|WOM��*C�����p�Cc+Uw��x]�Vޓ�/�3�&W"y�c���	-����
e�Gg[�x��6_��q߅,xϸ@��pr�s+�f����?��&�N��M��������F�(����Ӡ�k�mp�}&8��G���k)����w�����nEc\�")y�^�Y2 ��y�~��I�4���:El�PƖ��Y�Pu̞��F�0����Yc"���ZM��bqro�d7���e�L����7����Q�{�N*�NQ�*�+S�:=���U�䥁˰F�CaZ����p�"Ɓ/p�e��@����0�#5���C�ϒ�V33�:YDm��;l��.���C˖���q};�U"�*�0�d���;�55KH�OZ�~X�u�b�������T4��6����4-E�m��$�8�j�_��9�M#�V���¥�7�Zz�8zG������`M��&�e�|-_�55�63:�z$��ؚ�N$������a�oJ�����Oه��תz���ood�|4�q�>{68�W�A+{�OU�#�|�/(�#��r��P��o�R���ߏn�D��3�H}�9����۾Q	%dP�)�@D�m��s�^9g9t� y�/#�����Ԭ�t�գe����V�{�8�Gtb��۩���xQ5�3�˒;����q�����/�5���
�a{p��c���~C�7vv|0��7������Ե����=��K���"u\��z^9qķDW� G���I��1�Ω�pu����B[x���_�U���-��LZ��b�O`�Ā�q?�6��N]�"�#�b����+�)��5��P�^U�Z)dgrQ�x;�:�A�����rŷ�9�E�b�z����"��9+r��E��|���~>�P�t�v|S����%�.c\5TZm�PUK��? ��i�F�?�64��K�&���%)G��!��W-fH�7y7�%+K���m�g��a����L{��F�i|� _�Ս1P�ߢ;��]�b�և�1�<�9_P�&w��/4�n�vTZn1���H�Vkg�v� <'�8�r�ɑ�,���2儏
Ճb+��� �[�����"ZIqy�0�( ��`�DE]�ve'��1
���U�>���4&�{t౫���:��[�8��-���<z�Kނ!߃5�[�;�� ecjb0>�Vx}[���͛*�avf�l�{����4��'����K��侊��a����ڮ����q4����9�\be��\(ҥp�8r�V(��6�Ͷڪ98�M3`�<�?W�ۅ�-��%�O��B�2�)��R�%y��Y�wDb��*:�2"DB�`��@���n[U�����b~���$���R���g$�PΜ�6���ߵxՋ��(��P�Y��=������y�/
ΥC�!��
�m������!?�x �%�+�q��5��ɵ��n�*�$�P_Q������o��c����;
\�I���ci��B�j�p�'�s�<ֽ^y2��9?��ꄃ}Yڋ�X�Uj&�|���. 5��6+yc�A<�,��C u#M��E�Ќ��D��c��c�%�o�6	���f�}��\�SL!�W��L� �'G9�ȼ��9�H�*���a4~���K�Hl?,P���!�?�d����*������͸9�w.LK��"�,�x�v�<h#����=�tGX��E*�Y����}X����R�OB:JA��JԦ}:�eIv��>P�;�c���;ZIP�7�ߵ���_�;�V������p֎D�~�tM��o�3K��K�DZ��&�F��$�O����׾JK;�K[�|K��!I������ɇ䡠顕���tv�D�oC�&�\�}��ٯSOD�p�b��X=��� d������0�ˠ4� �uK �:U&�B'\~��kC���Q�GQ�o:e�A�
���Z{�&�0�e�iD�uu#�*���ћ8?Nx�[��$w��Mb&�ͭ�G��S9��*1����� ��nYc�<���#x�-�f�����ck���M�9Ġ��C��TΥ����E=U�񰩶��w�zՠ�6!�m�w:���d��������Utg�s�O�$h 4�ܮ�ʫ��5٭��6K݉Z�\|�:��T�fIŗk��#ىQ��iX ���	jĕ��#���K���w�g�����۾�s���`lc.��	��A�m{����1"B���rZT��z@��H��c�r,wdOQpA�a4H��+ּ�c��6��!���������!�'�=����1vgE ����<-����QNW�7��2w�E�#�y�i��m�ũ�v{}�n��SϹ���7�.ȩ�������6"��.��hh���[�O�rq��k��WF�C�56�RI�ӂA�m�w�s�l���w@�����a�
�P�����t�d�C�{@��$I�Oл��ȷg�ż֭O0�#b=�xyUD�����zI��F���_�p��/YTl3X�����ȝ���o��(3D�$�}<�[�*W/�	��(]��랎�c�K�H�ȑ9q�1����\�#ÃS_�|�|�����WL���
nTh�xDJX&�� ����I����D:��Ԡ���N����,�]�3��Z����2���R,�)�_�*��B�P����_�h��*;^9c.	��۝ʬ~'(����kW�Z�J-l�}t��:�K�n9G.���AS��3�"�$k�y�aG��0��:�z,@Tgn{><h�;Am*')�/�7ϸ�[Bgu�/����<m��~�� T���H�<	�j:��N�.铈�%���Q�q��功�Q'�v��m������Lù�dp�u4R�=�b�o�h��^g�/������p��0�bg��u���a;.��~��=@,�_�,�P5K�>�һYDS�e�N��x��x�'���L�*�}fE����	U5欄͐����u%k~5JZ�7�Y�bDcW�����X�#wDa0lѼ���knu��N�1g��e��C ��/o�<����,��`���Iy��-�\Ȫ��6"��!ݗ1�mSO��$_]���Z�´uM�(ɵy���D�?��ޠN��ԽRP\&A�CZH)OS�n�!���:Q(�X欔�3��H��%"S�Ldo�Q�D��{�Odgx���M�j�b�=�Gїu�b������"]Y��Ah=�����Nmq���2�������Fcʸ"LnoUu����u=L>��<�5#A}[X�H�ܫp-|*�dOF��Sy�����,�!���rq�{���3�H���E���4����#��L�}�v�y�������B��M��,c9��4%�8�33���.$38%H8)��;��lo�-��.[tk �	�3�Й�ڶ��p(�	�V!�	�Jn��4�k��w,n�m�6����ݒԦ��v��{���>�W�m}y˵I#�̖a�!�/E&��P��<�y� ��ie��cx8�զ6�k�s��b����F�3�8�l���m ���	��V��n݋�`�dJ��G��|v���c������b����-lP�δ�����.!�� �y��m�R�q)攏j�5�)�cj;��w�޵�J1����cŻCoI���ź$�C�@)$'�P^�S>j�}���v^*��[�L�a�ű����~s������^�6l!n��x�DC�
c��l	�j�2HH�K�s�WI�_Y�r�7��=/��(j�kL�qU��|����Ɣ���D��GC'?��߃�>e��%LϽ��3���o���?��.���˾���Ξ������I|�0���_�)I�ڀC2�i��T58n�x�����Qq�'����/�<���%2H�i �C���u��nd�9�9��|����e�_�+�|�wާ�MP֒w�X��v�if�BGS&Y÷xz��S��H���,�i�X�U����t�Ի�s�y��Ⱥ5D'��&�%��)��@�ұ�]q<	&���q� ��J+$8+Y;������oF�o�I��!����y�ѿ	���RC��/.o���RQt����i�5�g��[PK\��N���3ݨ����\H:X4��B�bEd����9?�D���NF���ǽ�2��b��A�C�zj��7 
5�ǐw�χ �S18J�x��v�C�dYP�t��֡�����[U�+M8j���)AM�mLNc?���(�q�u9f�z��$�-��'F�����Y�I��=�k��/y?�s�(���I���S��Լ�p��A�?F� �����!�G<2�Qpk8��#����6\x�-�FY��O�q9Ӝ�K��V��(�ϒ�b�q��i5�W�ř�BpDU��O��5E���E	�y
�@�%��S�d�AG��k��#�������u?F�H��ߣoN�߅�jTg�����J���e�F��ѹ��(Ye��m���qCZ�%���s�jp<\�?�O$<�$W�z��QJ�Â���=S��*����^����W�%Rl�N�c����f�0�ȁ;V�?�w��~p�l�t7=m���6�����84�'��!лtv�@m/�W�u�Ϋ6LsHo \{OL���ߺ B���b9!��y������0G(�-\�����88�|��V��qp��.'����.��8=���ed�?X�� ��7�o�#��y9�@��a�k&�̜8f�Z���W�����t�«��Q$�MV-��֗����D����Z�h���'[��]k��8����P:#�!�K'�+�Fh�{:��7���|��s��z=;��A�D��t�!���5M���= %������1��,�;ޢZ{��I������_qf��U�_���#�����$�0��#��){���'$�p�u\�Qd!W2���R��B	�h�v!��xEv����N��sA��F ��[�p5�]cv�]*�Uc����I�ϐ|���*'S~���U�b�L���?c=S���3-�`gN��\.���,phe�Z���x�t��q5xRS�	ݳ�b�)��I�.y;�u ���c�pz�R��p=#����إ��5>ɮ��x
z-�����L{�ҋ�+mG[���e0(� u<�x��N����68���Mʞ��{�Pu�e�������3xa#D �	tx^)��p��ؼBቅ��8�t &���O�1���ZxҕƎld���l����E����v#?	V�p����I�;�n����3<FS.���3:��_<;�N�9��N��R:Jiy|����~@���&���U���'X3|��̇�"P�ʠ]*N�\jӂ,���1�@�Z�"ه��M<�� c-���I�6���%K��)��Z^z+�=�ӊ+{6�c�*8
|��v~�0���K�͌W-lu�ۭ:��'ϓäV��MG|�����^�]�jGjf>ъ�&�:�(��л�w�}+G~�}:<<�\�U����v�A΃>��p�<��8q�QT��;n��(w���Zǽ>V���x�Z���t�A���N8�"��w���䴐KPN(���&Hhy�%��|�o$�)�x�P�#A�E��*��6ˠ	F���P�%��[�$l��� ��.Ջ����%[#�V>����K�l��h����Md��Ls5,4i�O��:��B�=�c�{�g|���D����t��6K���q3��R?�)��|�0A\��]�����Q�K�r�05ɇQ�8��RԮ1;m�yI���;�a�?�q�� ,b�3?׼���=����V�x��~l��%��l*1U�~Bc��sƉ��ݿ3Z�O�z[L3*0�A�l������vOsJ��Hyu��6o����?�]�b���?A̰h�>⃯X/�^��u�������Y��dv!:9ǭ��M����|�V�:j'����Ի��;Vc��`��!m�z`rcg�!�A�Ĳ�o�~*�u���~+H�_��S���Z= I��F)�1L������מQ��)��W�q�q��O5P��*F+���S�^Ln��$Cl2�e��s�
\������Ro8~(��K�n5f*�% P2��p�'&�C������E:*���N�.@̦]��i��,P�,�H��^���ܞO&H��G���H��	n����z�H`���~�Y����� �2&C�F����Bv9�K�ֵ�-!D2�U�#��^�V��|��6�X���`�E�Z;z�F2�>��7�b+ᴵ��,��ԑ�Qw:B�wɾdӨ�ze�{Z}^w ɑ���,�[��|��q��-�$�,���h�_1>����u%����E�6_}�\����?�ۘo��ivO��(� 6�1!����Y�����\����@�L����ma)_"�X�\�
��8d1X��CT��V��ڤ=��:����`�>P*ދ���U����j���%v5�o�\��S�	^�&�Ko1ƥQT�w��m���+=Ǵ�C/��������?�����X�F��7y��C���W�tW �7�NfU�<ojk/�u\�U��E*�ߒՁRg�������*1V�a���X�^@(vv�r���I�αR�Cc�s��4��N�?;�@���{rO��(\��F�q%� k:�R�0�N-��
���c�����*�sMTK2p�{����i�� ͕��t�-���	eT�}
#ƺ*L�&?r�����(�0 L2 c`�|7ų�,�J��حb����'����g�Si��	X�7)������M�@#�M�b��Ew|���)���[дp�)�lSI)��=AAl��ȔD��/����zo��"y_6r3���7ޚ(��C@?�6���j#ٴc'���:��+X�
Hk�r��5�E���r؝<�
?�H{��ߎ8xk=�v�>q%[����&`�~z�a0,�?�qu�MV�#��nW�����P'^U�Q6.(&줸���c���S<�y���%T�����tZe�K/��&�m�2�P2ߞ5й�ipgZ����'+I�l  ƞ��h�^d�,��*��V��S�!���p%����v,']��&A�b�s)a��Ҏc���5Y��n$��t��Ce֪��)u�x"yh�����At��2K��h�`	PiJ�*���f�n���/��r{0�k�ޘ�T�o�q{;%���������?J ä$�S �fɶS! �^1T��Z�`�q~���3{�
u�ֲ�O������./��'�sƙ�(<�3��lGV� "����I�X�ՐhT&j�kT^��1Ŷ�W�Ļ���~��8�3=�v<)��=0����xs���˳|d��[w�
����e�2��4�����
=���@�$�����.�=�+�p�5�`"�;/رB��j����|�+��ӈu���:��?Q���*^5��kc��3I��䘘�H�m��/�Q�j�s����?��J��.VD
�!��h��t����-yX�>�+�9�̔h?M�3�d,��'1������03<���Y�u��[u�r�F�����z��X��j��Y#_�� ���T��.�!\^�W�ůד�4G�UH�-_���CG��}�IM�ʈ�����2��
��d�7D06vR�Bm
Gؼ���T@�D�q��hV1�yA��̱�:55�[T�c��!~���h+��老�3���������T0�AW��Tq���M8�� ��I˖�;vA��ǳ�]&�~\�N}=����Yj��H�!g��h�)��?b_�J�y�H��I�y�΄�H�d��#u	�|q���8�:��9�!���\$��<z��QQk>1���!z����+J�rFJ���=h�3kS�t�R�q��9a�I��tr�}��t*�M�+���Tμjf�&/�
�ڞ`��/�!������=�Įj�jC�gWL��\)u�0�"����%��4�W��{��sp�Ͳ�&^�3�����?���S�l��?����A�am@
v���hi�ܥr����,�ErCX��x=�?̆h0>E�Y�FB�wf������B�H�ەh���E� ����8���	嚪�ᕧ���\/����rߛ�a����|���-8�EP�sͭI �!6�M��,�A�
tx��wD�4	�;w[*p�c��f���E����-��`ϰ�D}�덣W�C�����ɏ��} �o�r�I�����m����ԇ9f�"F�p[:�\"�Ё��.�V�����}��B)�m���cc�%���x����������)J"	�dx���쐞��5F�?G~��=Xt,(O��H~.�M�����$�j�dA�4���5����ː���O�J�3���^�mue��:~k����KM��X��~�ן�H��s(/c)��Mx�QS:� �R���Nv4GYh��o^���-���@�XyYYA�vÿz���T�z�L�U��Ȧt��(d�����BП�q�f[?=���BgL���b��w���*e��-b��r-��hf�(Î��g��Y:eP����0��N�x����Aʟ�3��g�3f�$��oW���PG����� d���i���m���1�������^�9��Z������iNgH����:)�e�Nc���U����D�}
���2~�^��?��c�$\}�h�(2�C�2���8��1���J�7U�?�V�R�tB
V����9�g�ʢ���?ڻL䇸[�R��\��S~4�3�m���W�i_��qĦ�7&n��XsՆTPm�cR���Qӱ��\�P���\����<Vڀ���d9������N3��n�Z(is��΁j�b@��v5���n%)a��*��4[���l�8 \`s�z�۩C�Kx�S�N�����f+���-��6Ϲ������L�P�ɮ����+[U	G������gr�'���Z6��N.	B��sڈ��K����"���x�\(�	��ٖ~��pԭ۔��s,�ʡG�R��=���?Q��: �W���x��d��/���ey�4b�oH���扡��a2��',�ˎ.�mSӎ)B$��ȕ�*���Q<Ǿ�"*ʟ}�\ߙl�MيS[�M�L:���M�ԁ��/��@����׾)�dL	����܈����u�\��G'wK�B�'�1)��k�p�{�r�N��s������c�Y�'�KR��&�)H�4��bb�YO���c��Fl��G�O����(�k��� E$*�f�sY��� /f.�;,�8�q��iW�����6�e�c�)5���R�ӗM��%&�C����=*��:�_�]G��0=��Uq@�c�z̉ ���S#aW�4�i��x��=��y�I��X�1q>�?�,:;1Ǩ�,��x��'v�GTб�i};����Ei��ߩJ+!��m]`[s��K�;ȫ�M�P����+x�򢿕�(��h �(�X�A��3N�I���%���B��ǿ��j*>H?�#!L��J;�DoeAl������C���w��+y����'m�وT�	g��+3Ȳ@� �O��é%Z�lś�����0�����*���զG����?�V�1ر	��  B��ƅ�;P#6��ի��9k2h��TYe�_b�s��@��[���d����yG��q���%Y�"��^J�M� &9ez�l�x,ɥ��S���.ږ�bKn�ܳm���=䃌�S��?)�*�Ra���ӢR��M�o��֛���z�l�,�m���S�ŷ?��5���4J58�Q	'����^;L�}�@Y��%�ah���`t�\�zS��M�YZ#�����B�]
/Z�&2�4��(�+'}�ޤ����~~�'������d�:��xd�d <�y���)o�N��ek ��B3���aa��`���_N!�mTt�6�����b��y�O�=Y�I�����EP��o�TD����e�C;vS��D�B3I,u�����Q�<qB��.���Y�
>�U�K�jAY�hg&�x��	���a�T�;a���@�/��<9�b�3_�	�a�̡Π�ܚ.m@E�Y��
� �D�;��R��릢�$�ޓ& �<q�:��VYx���y~��Y}:�t@a����j�������Q0��/r���f6�.��K�L�,��ܚ#��_���S�k�w��ˮPbyYy��VGX{�|��5N�j>�`�_���6�Y���6����Ol��
�NY7�.�Vm��/�x��W���<�&f�p�A��1�4�E��u?>�������M�k;�x�ū�GJ'��0F�6cn9U60��1�@�d(����V�����/��%]�2��� 4��^�~��d011���"P�5'l� }R!E���`���'�����ct�X���v(��T�:P�D����5Y�p�DO~SJ%G�e|�o����&)�,uA!�h)��z�L|���gô5�����k��b��(#�Pdl[�i3��њ,㑗*��:��j\N�/����»���¾y���A� N�
:׏����1����h?�%�#��Y�5 xP�+�Z������\���9�w0#+�p�l�(]|��^;9D��l'm)˰��wĜ�sV���P�A�ܣ�u��]�?_��q�qAE���+�XF�Uwe��izyV'lÃ�x��^���������Y��K]����E�рp�w�Y{(g�ThzY�к~�K3XC����ǘ�MS�uS����>ǃIjVF��@uI=��Q�o�Yx:88}��KoDSƪ��1�y�m�n_ļΠ��<��G���ٺ��	�ƞ�L�Up -%E���Tϥ����A�>A���[���_�Rr��"=wi;��K���KFx�ٺ�ʊt��r0���r�[��Z!������w�>�RN��X�Y�x;�
�7��ᆲ<��$�`��h������,�E�챱��4U�ʅ,�~?��m����#6ԴzgFIZ�1� *���G�{�l�#���F�.^i�!]�f���`K�7WE2��YM�젻�����1ₕ,��l��Z*ʷQ����(:*��!)Lj��Yb��ӹI���
:S���
j���r��T�qN�]gw=g��E��a��-�.?���PR�*�&,ۄ�W�pb@	��R�Ƣl<���e��=9v3ס�?|l�l�Y�3(�d�ɍ���w�<[؇��UaX�x,l<�"���fQ�40��D	��rơ�[��#� �6�R2euW`��{4�8z��K�B�i�c�����`ϣ�IЙ�f��݌�n�S+�>�*Z�{���CN"B����'��R��s�fĿ8���.��A�7�}u��dg@�9����I� 姊T����e�6�a�u��7�G�	s�9w������k>Q�g�C�řV�i?��U�S���A4,:R-���^'ߥ����}22�^Qzjߑ�{��=�����m��._��`V�6DF��RHEqR�� �n`��htj�����S13��'G�BN����0���Sm���K[��a��B��^�1%�.�	ȗ��W&*����ۅM�[H�'o.T�x��1P�j��Ѕ�P�gċ3�%9Y�KLuܦ������>sT"�H�Du-�}�d�)�%�}���o߉ ��i�x���e�7S�Fm�pЦ�7j˸����r3oH� W�T���"�*��r�8,�yԯ����A�W�]���Q�.��/m�h��h�>U�G�)�<8�����D��w�x�u�;�{���X_zC�k��S��6��$W���wHD�\o��8����cb���?Ҫ�F��U�E�۸�oh��6������@+Yd��D5�V�a�i��Z�Q�+Z�Uh�����wg�|��|
��?�1�}	�aw6~��:vL�/55!~�!by�D��=��ړ�;S�]��:x��F���w:Qe��O��{6����[R�S�=gH��F�9��.�f�1�r�+�z��(�)}�:����t�ˁ��K2l�5z*���z+�<"�lY���dnh�l���YL9µ��\m�
g��
`��2Xm�D��C�y���9�_Q��7�yGi�����?���;�R�j��(̉X�qhiA۰y�XI�W��K��Kx���Lpo��å��B A� �?�i�V�v��b�[�� g��2�l�m���ޯ�?1Bs@��Z�.,2�<}�Æ�pA�=�[�E��ܚN�DXuW�7>D'�Q2�Ac#��r}���7�U��p5
`�#"`�$D`���[9Ǫv�4U��t�PA?ݡ�,������$���s���o�{�V2���5r����u����i�B�t �n��~�DSq�<V��mҋ�ׇ�w�3ݾ�V���\��]�W�8�����f&���	��́g�����T�R��}+m�o&���1�\v׎Nt'Lr�[w�����t�ۗ���q8�w�O�>�)�z����TPD�+����BsO-Y(�z�3���g)}vW��o'�.�`{�����`?9�`!�G�N���4im]4��&^23<���'RZ�M�Hu���s�`.ݽw�)��$t`�q��Bw�5b�́�-�V���%h���&��|2Jg�*':��*�����@ �4L�CQ�Eb C��H���5Q$����"u=�	p�d�9��t�C�oX����WI̔ĄZc�xb���>a�&��Bx�t���b��kg���[�3$(��4��.��t��I�����Wj*�=_|�X�O~?�Y�x��Br��^��c.��9�ّ��y=Ade7��B���y0�� �ȹE��9�n̓^�џD��q���f@���|̧A�o�
��3tJ�u`�D�Q6Te����X�؞�p�����4-)r-2�o�cG ����d�`O���hr����k݁%�a�Փ�f�4ʝ�:�6;�Z�nYl�H���f���Px̚qy�\��^��
{���(xx&o�4�`Q�ɞ���ޕk���Y�����aΞ�� ��q���?��;P	��F""�%g��4�	EL>H�R���*��xF�(r�@�M zS��,��C���߅y!���_6!܏wG2T��R#���V b�dr,-�S�Z`78�r\�������O�	�%���n�N$����f�O=�0;������1ӝ�5��Y�*@	�y�Qs�Q����7�Y��).�=�����a�eW(�G@9����xb�Ǫ�c�Q*����;CK�f�"��9�����D�8�/���)��߫x[�I�e�a��>�����l��$���>n�Z,7�l���f���0�.f8�ޞPIc̈́�2�th%C�g&��s���D�kii�snN#N��jzA�/�z�'=	
�;�1X���cn�l'��#C+�#��$mBnWB�*�T�!�'�B[��{y^���<�7��.̷,��)�.��E�<�������n����E�D���_8G,J���c��.�� |�DƉF�]^��f %3*�#0���7R&6H���)"�[�c�{�r�H��&�P[M���P+�����`��{:	K���,�M��ȴʾT[��:�e_F|�|�Q�������B�$E��ZӬKˈ�'/?�wөYv��5�)+���k$_G����ЪO�WL�)��Z�\��+[b��ڊ?��~��kV˥\�n)C���Hi[�j�j"N~�ͭD�(G��ť[�4O՟�45�,Ρ*���}�	§�8H�n��{X�5���=/@B�ۄΙR$��[�0���x���g�;֓�B3Y��ft�(rC���Ui�8�2G2����پ�����q/�('U���Ḧ́�����1�n�p+��+��/�c��±��7N�m#%%9��8���U��.0\T���)m�] >b�j��G �U/�ȏ���W���K=�u�w�è����5/Q�;�8�����q� �%�he�5� ����ن���e8Jg�PU�ȉ-ZʲT�����\
	�y�n�kk���j�9���F�o���$82嶔/|�8le
����G~Vt�f�}N'���rK�,w�G�%��;��� �h��
zH�o����}li��� ���-ej���Ԟ�{g`��nl�u-�23�V�pǗ�7�Yv�{kr�w%�E�2-1�\�^ơ�Ji��� ]*&a�~$L��\����TTm�X�Y�&�Y����a/��GO>;�Ǹ\PB���=���z�LzT)i��d��
*�-a�JU{��V�TK�P�}Fa���
������e;�/UT�ɹ��qe_��F!wр%�ؘ_�����#A��cWZ�d,x��/��4�.c۔�oT1V��-毾�H̉5�4���E��5��X��S�	�'笂S��i�a�!z#���UN���Ƙ��&. g��߳���#�jPp0�o4� |��T�y��z�Y=�s�뛬Ďv��ήX�HW(�?���0�Ϲ�LNk�Y)APZnl3�	?�=g��୪+٧���Ѕ�v�'�p�~�D��J4�p]��_츎s�i�C:�(��&�&����O&DǊ"@�?k�������l�̋E����XѰ��;ϫ�¨w
�cE�5����à�< gL���z;k�,���ʚ=YDՕ�U�9��]g ���[L����[��x��X��B�La�;��K��'B�B�s���px|�����R��j�!�9'Q�_�\�~ ��Kq@Z�vm�Θ'��#5+M·o=_[hȻU{����*s��U\�mQ�3��!��n�{C�ZE�Y1���yg��$7��,ܓL�bD�m���eӳ�5�ĕ�����N.^��'�Ds����I���}���b�M$e�>�6&N�E�X�P�]�H
T��$v��sM�!��؂�X-���|ߨ&��E�@ �.��'�f�A�o[�f�y]"� �d\WT�i��U��?��5�t���jK�5��$�#8��?�G����wXgǭ��wF)���FJݶ� iJ��3!�yJŏ�;�G�j��%�FU��Y-� �����@Ӓ�x�}�H�7Uȉ!sl���P閝M�s�,��U����_0�t��P���0����[�K�o�i�6K�h��°	�H��y`w2��G@��� �H{��R�ӛN���i"��ԉ
V�
�
����x@j��q]LT]H;�؍�.na␓���i
bD�������:16����փ���n3[��eYcS@0��U��r�ݏd2��׭c!	�!l���[kE�/W ��a'Y�W͗�UW��D��t_dpؼ�7�~(��7�4���v���}��沉�d��T�[�sb���
VZ&H�<�5���g�y��;;��c�b�e��łcƐ�4�� ���5�?�{��ּ}���_��T2ן���n!��a{���K��	Y��<���I�eO�����!��q�2����͞��$�97�U}��c�)GFRE�J23@�21�4>�K�6��vt�{��"�@�J�ݹ;����m�8t�"�a�F��*��ԓ{(�F���W�A�����[�P���O�T+��&�#�4K�Z�a�5ų�VF`��B7��@�R�zW ���;�	,���������q0����J�;�X3-�&|�E��`�!�~ʩEADXյv�J��~E>�J�tTH8����I���ZO�+�z�5���|���D]ߤ���XU��	��b�\�D��TV�ZצO����D����3g�{Z�z:���V� }|����.���<W;��a׵�ij&O��VϜK�������t?lQ��Ǻ�uި=Ei����m�e~��Y�L�	QwK̝͢�Uׅܲڰ*2��Jp����R~��i9'e���,ua������Y�ڮƸ&e*�#�ǴDĿ��X~v�@�O>�V����KY�x%<*0h�+�F�gۤ;���#�RR��xR9 ��q56<{aL`��4�w��2��J�ީ��G�/����q���u��i���g5���6��5L=S����iV�(L�Y�T�DC�����%@�%f.��}��>�x2<�����K���Q��ş�1ۇ�_.��y�
Ix���AD�5@O%2�5z���nK#hp�r�ݟ?�ޝ�Ύ{�x�%�t%Έ�������H��1����U=0,����(����2�.#��Ǚ�����,����[���O��Aܧ������ fJO}��s�#��vi����A$��Y�� �0ڟ,����7�n�JBԂ]po�+��IJF�ﯸ�^\<[�"2!.�>H�AP��x>lKi��6�R5��?���_%�4�EgY���U�{�x�u�}�7*tSː� �����X�KU�w`4�u����Qv	�i��_W!E��n`�+_uUG��uZ��Lhk���K��C3��c"��s�/�	����z��/i��K[ƿ�o�y�x�Ψ�3��cXLӑn�#��7�%��'��r�	v�;E���2Zzr+���"��7{�3j����;۵N�X�lz5H���yH�i�S��P1�V�z5�%"6: �=����.ER��`z<��ܭ)ڀ�_��dQY!���s*���i�l^]�q�p�89F���Y+K�i9�,�a�F� Q(ț����1�2�9�D�[��s@��+�U�������v�e���9��3�)�^ �c-b@��K�*���,��-~����Ů$��CU�Y��zg�tq���1<���6���C�K�K�+@ι"�;5�F$�]�:���� d4}��3�V��F�2[���cB�wG�i0�>	V7\�2:�L���G�/>2HK���xN+�*G��T;C��V���"s9�����4��	д��RU�Gެ�<\�t���7�Q�>Bf;�%�Q���o�8�&�0xPc��mHN*��6P��@CՍ����J[��ؘ���*[�V:;O[�@��\=[�����1�������y�7�Nq�Xb$�2]P`~��Ы03��0������4���(��Ւ���E��ž���"*����~��\���O�2��g���z�Bc�ˏ	i���)EcT��!l�h��z�Ҕ�o�8�Kϒ�����x�ڰ��0�C�t��g5��Q�[Zɲ�#�hN��a���c"��p\�^ݙ��׆�H�:��<�l��QM�)�x�ML_������ob�Ҟ!�TfX[N��Pf���y>�ȳ_�q����
ͷ�`{�ہ�x��B��𥏽X��Z?`R�����?�j� >|��*�9��1s�.�.(�k���3��C�y*3"��
������&�MO]�_�g_|X�X}De�ݝ���#�qi t��v������S�c#���3>���W/2�w�8� +?���@�~<��n�ܯc��ǿ���C�_�������@�s��Z�x��{�Ƒ�gc
�5�`Z��T�T�o�EjrUElDkeoʱ8]�QY?�%����YC�sN�l��.����r�|J��5zZ~{�Vi*����VFړ����k@?����4�4�A�Y��꒻���=�f>��`�>њ=�����҇�<KV������H�}����W(������ޡ��"k-�Yͧ����k�HC�D�a{I��ٱS��i��m�b�+�J98�""��Z�����*�D`F��6q'+�����n��?_	���Y#Br��r)yaچ�u��N�l�2��G ��]��8I`��x���OL^���OD�r���*���$�v4��2��������I3�c��ʔ��/�?#�����?���s�O�s��mF���]�|��Z�70b˜�ʺ#5�}�h�`"����W���@��I�u����hĴ�S��x^?D���{E�ꕥV�NnZ���A�-_�ũ���L*��?�!#����v��Qʹ��G�J�/�⎟����3��	�a��:����fM�/�b}5}*-��a<=K�^^9�	�M�D������*Lo~lD'��wb��c�k� ��!]\�J+����ᕉ��<F��ܢ��f0�9�����L\]d�=;uo���	�}�(����)?߁<�R��x���jM#��P��
W9�5v
i��S�r1H0c�[C���f$շ=}�T�tH:��eٝ�P�[�6o�w{�[Yh�Q�i:�n����v��F�����S������\��l�7��"����$H���ķ��(���j��K�yDo8���o��Vr;����?�	X~�c���P���%F��\���အ�����qZ� Is��Y�:+�����L�+�/B]s�K��e�)fZ�S���W�ޔ�4�^9�ęD�͆�Soס��z�~@��$�ܨ��&���Q�N�����1~�(7�\XS^�	M�4����H�=��nq��r^�内�ףːjGQ�X���6nu��~�Z4�!����$��9�Y���H���a�!��=�&Tk��n�� TR%S�O�����Z�~դ��7Bmq�]�DqB�G�=�}���`b�D��4"'X�0�2�bMY^�Y��Q���M�h�:P�r���~Q񨙖OCQ�Ð�B_O_��Yv����P~���s��j"I�%x��w��Z�`��W��j���n'� (F���D;h!��©���Տ'�>I���R�ԭ o_|Q�������ɚ݃E�]���,�
?>
������Z4=��Dd&�xp{s��O&��pz�+�� �� ������5i�y�U�r]Rg��(����E�,��tJ�V��YI�9��L�R��.�`x��)�T�sP ;��X��)
1E��Ԃ.h����u.ԋ3��i�XbN��)8��X(/�&�U^�b�M���� E��TO�����2��
�6���5XS�|�п�6���!�mp�Q���Ƭ�S�Nt�]���Ĩ~7B�{��5\f���� c ��F��u�N�G=G�8b/[h%�"se:��a��H�bf}צ�O_<vLZ���������;�ͤ��68}�X������8Ww:,2��6�8'"~�����;�{�H���U"aJ1���b%��]w6�k��3���FT�`�'��֫!�����<���i[��G2�Ƙ�T%� X��kbU���rlĈi�Bѩ���+@�?�R����%\�xH
��>�}�7Q�}�&��x���~�9i��0)�w5�ܛ�����פ�^ޏ?--���&����vc���`�f^��B�g��~h��L!��B���ӈۑ�6vUA�l��M������L\C�A��2��m2	iQ�#�Wk:}�|Bg�.*��q#`E�V�qw�K���-�K/0A96�V�N�T����U��~~l�*E{�Q�3�~�NF\�e�ꎸ<���mL���� x�3~�T[,"#�ߺM�q���j�`/��oLA��r��eg��Uy�)͆�ܓ�Y��J�C1 �Z���<��%jy��r�HW���(щ�B
�X�~�Cb���Xf�;�2��HA�K�xFe�g�$���m*絊�pT`̉�2::j�':�p��z[o[�
�$��P)Ʌ�'�,�q�Qf�K��@�p5��!1��W�vB����ڷ�l�ŶTJ����6��f��AU��Y��4���G�s�N��yd�� �0l
w���7Y,&C� �8qw���\1_]����*�B?��h���d�^>M�g8���V�ؠ�]OB��U����pM5�zh�A��h����.I�[�zڵ>o���F� 5GJܑ���d_�C ��cUD0�=�͢:OU�G���`����� ����=Ua�|w�r�Æ�,�A��1Ħ��9�9=���Q���2��D�k�n(E�}��n�*��/0n�gr+r�^�]���E��1�d��c�[J���)/�����졓|���G����`�6�b?Ȭ��ٟU&�u#��Р���L�%/P�g/T۫s���"�܈��C@f�e8�#!��I�Y����O��@�������� ��}P��eG�=�<Ke,�Ĥ�e<�[zF���1�|��騬]�.��mk�WO�;.��(t!�\-%1g�;��tn���o|fnD���q_p�z��_�n���0�"6v�C; ���Ł'�t��W�[ܷ/\,$�vR��@��=����l��� ���y�<���Π��*�ht������]'b�����n�Nd(����B��(���k[p��q��y9qz9�jLX�c��@͕`	��,|��:���<����α8O�5�!6����h�_�a��=0i�y�3��a�剳�Vr]��O��&����\Rc!_���N�F�B'�[y�L��A�x?��|V�t$h8����>�E�����O�L�Z�T ��ܡ	�v��S��gB䥻����,�\��`q��:���lO�/����J~�'ڳ����Y忊\��x���Je	��8����&��m$�KDO���Web�����~m����B��{0N�&��ϻ��?�Vr�,QV�
��pP7�D܋�RR��t�������7G�:�-Y�,��븜�ӳ�1�����f�ed��r���4c@C-�����M��B��_�%�Ȝ���̊Pm����XEF��Ɩz�����n�l���#C�#1��[� ;��o��*�t�Ch<ݭ�<�+�|,�������
wT7���؞�"�ތK_�&��ZOG��:�՞����CȂqs$�E1-b$k����tTSp��l�VN�`�R[��<լ���6��h��IkO=P.f�y��K7�Ŋ\��� 5�7n�����]�&�AZ���{�Ӄ��1~�-O�˼�ǀe�TK�@���'��G����M��ʿu������4c=\�;f%�3��ȳx�=�)GE�W��v$�Md���g�ȫ[��R���ι~�[+��W�7��u����f07��0_֦su�MJ�b�K�.w��FG���� ��xfDB�����b��ę�� �V����E���/F�,�U�5ks�/��R*vw�xB����\�1����R�h4O����$,{�D2��s=���+�� D�bi$�
[�Ŕ��B~�҇���;M�zb;c���r+��o3+�	�>�K�����0��}�oqf,�������E(s_�a��/��qG�1��=j\������mU���<��ZN�ԇ1  ���'�YKT��4�de���@K��>~C�2�0����	�"��"��X�h����)��޽k^���#�I��b(���ꆙF�������v�m��Zlw������:���/4�C�F,5��F�PAۇ
g� �7Z�"#���j�>e�v�lZw\xI��!��#�����^h�#Ү�;�m����Ǐ��p&�TN���{�T�qe�֠��b�Y�t6�S3[U�#kZ�>3C�0Q+�k��Z��`��6���k}�PD���u&���1��F��fR{�5\ʪ:0"����cר�"
�(�M��.�헍���N���9�_8	�;p�nm��D�K���2ٽ�V�A]RN��Ã�j����S�z�n��س<W��vS��d}���h�{���;*k��U�R��8;o��:P�)�4F�/�sB���Y�:6���/�i�ΰ�h&��s�r��^]�F\.�@�BG!�/ ��Y�����������;�>+p�p�r�����i�Y�%�ɖ4hR�K6Ս��`�sn�~�Λ��β�����؎��! �]�0Kv�㢠S��{H"��nM��<Y���'.������b�P�L��$�K�e�+����{|\�;��"���|��l�֤����&�.�ܓ�2��p5��H����@ �֕x�3��⾥|�Ey��O����$�j��q�oPIli�׻mtb}������v�B�칗=|��W^�,��^zO�Y�	���}�a��b5�4QG���d����A�&�u�RS� 1�凼��ኪ���c�1a�+]t��
z9�}�f�'���D�A�ƺ�`t�3Pz�3+fa ���)���yKTz�Yn����9j�E�i�����/�`̫�jd�Z{g�I�%�p@	\�rV�x:�,�"	DY%��FcK�F�)�H����~' �
��1�
$UMqߧQg�� ����c� Y.�I����g^0=C����RR]p�=�[9�|O`��RL t�zm��1R�Z�w��^��p�TǶ��#�� 8��n�=��B�nz�d�Or|[��v��!�9��w�خ��Cmy�fА�	�h�3g;eE*���c}���Eܽ�Lr�9�z^&�[�{[��af��.U�7�=(W[�޽b#46X��ڐBC�瑴Y}� ��P���s� W���^�G�|ƞ��%F��TGϛ&��"��^���}մ���v���J�_�����*4����_0��<�%�_�Li��>��j�G��󷩪�8��|��S�Y"Pu�*�%��s#Rֲވ��'"�eL3����{�G1Mu���YW���x�?Ц���?����l+���/���ì�YE��G�W�ͣ�F�!�4_��YGc��Kꎣ|s�9��w��$-��Lu��uc��;�y�Ê��Gv�KAh/�����`�/Ǩ�����t_6�m��j��%�2�**��#����sAF �q��=2�R�ޭ��Y�=����h�Π��<1Q�P� N�M��h�VW��a耷(x����Ȃo�2��ѳ8�f�p�A�%�ct��Zt]��
?��K� �c,�C��.�=� ���$��w��a{J��@Z�|�
��I���8��W5+O����٧Mvĭ Q��V�&���v�C�����f�g"���	`��V�ΐ����9����/����gT�B�ILfnNB�hf��d��b�E��	8F�6���u���7rW̖t�U����Q��Mtz�f84s����r��xp�zcH�+Vk-��x*���۫���~���%Ɇ�Sv�������C�hֿ$ɫ���6kk5y&�`(��b�+H�"x���(FO�� �t��:�Ck�z��H4����ˍ#�JĖ����\��CRDmg���YEsiw�$��pS��$ba��`�&(�=lO�(h�5<cbҠي����4δᡠ����)�(��Rli{˭�v�ͻ�q}�^.D����y#���d�͡e-6���]���a[?��o��#Q�d�\l��-D}�Y�S� ��H�ɂ�w\n+̀���g}��z�@��ȃܤj���W��v��u5����$}�.�sK�D��4�����o��盐dﰶ@K�0rzc��x��:�]�����#�wt!��EH�уy�ĈU�݇��#��eǵBa�J�	՗��v�g� �̹4�b��0BZ+��e@�9閷u����[{S���}���ZƊ��0��궖��5����V�EXD�ዔH~�~����X��wxYь�%��y ���4�=
�n_��VJ����+��,�c�*�_���4T�k�=���p�|�_!Cl��M�m6\ O�" )�d	�a�v��k������N��^O!(����L��ht8�j�V_��p�R�S�� c��Eqq��h���e��0�����"����K9��Rq���J�9�Ek!]�aL���r�2���y�j�� �Z���rF���!@z��A��DF2�7H;^�vh�0�F	$&U�I��|�eȯvҒ��*�T��߲�������6����&I]pk�8V�wT�N�Q]F�����|���j��8�_���ͧV���\I����.���1EU��Rg&�`��6�yn�ӊFBC��
�t@"���J}/�)��Z�V��"+��a��Y�FTt<)H�e��m|�r�]��i���FR��ѿ�x�9#K���
��7��E���웴��1�f�Xs�§~�&QE+�`�Qk��I���pӧg�N�Úz��a��4�v����I����/n.���5�s&tiП�G�Eٶ�-�&���E����j��Fb���6{p�j�d�B
�U�0Qa�Y��b�N�UÇq�0	()����|��F��"��&����5�]�/H!�X�|w�Mh^���r��ع�kl8�*�wN#�N�O�ZS�u�utטTKݗ�;sjC�]�;�;�[ ��N����;��͈�=�FTpJFY�d�Ӎ$  @g���QVK��\��R�a��jH�1���큖I�?�v��	��%�՞��N�'�AQ�"����T�
�����]�r���wP�q��]+�K4�����B�E��X�o��_I�Α�J��%�wj=[Dm�L�l)�H�0�M^��e��ߓ%��e��Aǅ��f=�aayÜ��-����a�'�y�RBO�wC��<�/������YmDzV�4��^�������l��#�%�S~�xB�W�8uU�Be�X t�ZZf��J��ݦh�d�߀����o��H+7떷��n���x��W_�᤹������o�Q0nM7��������*�Td�B����v��%l�E�,��`�������1��.���"S�Hm�C�THOC��lR�����[��L�%S�Ȩ]~s���C�y���������g���j�/8H�I�n�Y����4�6{��y�����l$5�Z�)�z�|,Q-׿���������	*���n�/�$w�a}>?�U`���F]�% � ��=�Ə�?��i�)��/i@oV�r`�� ��K����{{�*�6�����o�sXtJ�5���H�}��6��#��jȱ���/��,����[��1z�2c���q��ƍ��4��n�v��z��>3��YU�2!'�h�y��V��WѠN��
X�1ɽ�Ib�����Ҕ�q���fX�r�)�AMCS,�N�8]b��n�XЖ��F@�w��	�qC�W:b�:��ԡ?ޣ&6�����j'L���~����|�į�ڥ�N��:.?t|�@�|�?��CJ���*cKcz[���<����c�����Vw��1�|@�P�7$��<�}\�yBv��e��YjPJJ�ʩ�Gg˺6(��4V������q�I���	����6}��a(��5����6p;����i�C����Y��D���$�pyN$�����eC��m	z9A;Ly%C:�B���h�:��V����4d�d ��~��ZvT�W��n.3�7m�I׵D��b?��Q?��1Ecm��$���1�ݫ~3z_��a�p��ʬ�Ox�7���Tr�^�����F�FRJF'�~'�'��'0�ڣ����z"Ò�����7�~	�'�3�;��:���Mz�M�|���[J�;*W_�1rr��P��S:�j��gI�'�U�P�1Z�9r��
�"N��s��k�	����("n�������T%���"�|�O�p�A&ÿ2��xӣ�dv�^-"9�bF=�#s�e_�e*E�v�Z3S�M�ݹfd(�u@s�\��t�n�"Z�����d8���
�2��g�_*�f��5�`Ͳg�Q?��i6i)c���luO�e��P�u܏�!X�b��u�/�~3���ވ��0FɎ�E����b�~��DME|y�c#ﺉfǥs��3��l�P�0at��F�Z2�b�&�f���J-�����(��&v�|U'c�����Ib�*�m�$N��*���OU�P⟥B�<�eG�82'�\J����&5����K{Ŗ��/������4��n�݄^ś�z@�3�pZb|�@X�N� s���T��x��I{�g���,�Ň��˳}@5z/��R��VnB�+�������B,��/xO
C|u*��CŶ��k��+#{�J���y��$��9�1j��M�����";}s�(����� 6R�.3j�w���)���(?��2�aF\�#C����i6�M��q&��<�u�qkGOƁ�!�Jfw<Z���z��F��+�7䐅,
���X�x��H��=���F�r���=�� _d��'t���!YC�F/��;�ld�m�w"����@"�D��d߭�.�wWe�`I���� �����Gm��{��FW.4�Q�2��]�c�s_h�(��6�0�,Tr	i���2]s{֯�fRui ���.�������c��"̪- ���mWP��G��)�B�3'�m��LO����a3���c�3$ DXG�b0y�ѿQ�n��kQ�a����.�*8 �C��b�XO'��,�'u���P�Q0>���M�޶�K�4�	z�S[��X�1�;ד��gSP�*;�:��"Ӑ�8��ăsx���� ��I��>���.tG���t�G�ү�Ak4$iK�x�A��W��L9f�rhu�v��	�N��:�U㡖X�?>�D�H��p��K�N5a��R3����s7�e�߬��6T2�ɫN�%͊?����8��!v�Ŧ���ᩎfҬ���\{��Y���d5��"A�O��8�ٍ�|ل�[y��4G��
4�%�d�'�ͣ'���<������P~C�Y�.n2|�	�E�gˊ@d7s���<����ŷ�Z�`���2p/0����(H��5!v�,.ii���q�����h=�nґ��'�GM*�0S,��������c5�U҉6T���5�F�2��pb_ǵ��I,����zlոd~���|l��.$����iⷼ#��9��Q���5E|PY��Z�G�������"�칟�� N{b����{'�c��ݷ4�k�6��� � "�.H�y�]��Lb�LE����uW��LV�I	��'j�{ᑏ���n����Cy�;̡�H��]���t"��y��＾|��a����}��#���56.Ԧ�����%�����$��2V��`�^)Ka�����U�&]s�p��d���-̓B8�9/4�@��p	��B��.�B�
���ǯ�)=��x�7b�n�z?�hX�ж��:N�9 x �{c��#��
_��+�lh9Ơ�g��Yv�&�M	7zP��7�dupeɻ=TvRD����^(h��_~��ލ����40���5�q��Iu�� X�p ��N��x�%g�P�O@�P���R�,q�qA<���s�����Sr��G`�l����g<���TVGR�I��]Q�]��ܻ�n�ac��dXJںߖSu�B��%�e�Q��n�U�-$����ɦ��Ļ�S	�G����|��J�|��J���@z�iz���p=�ؤh�*"��/�tbD�-!�ѦdW7F����gYP<WJD¹���m�,l�n��1�,�2�!ص!N�C��@	+n}������"��M�vl
X�`���8\�:�J�(�j�Nuj�q�\F��`���G(&̹l��J��DƬ���T��n��Y8B��ߙ�������}��?%4�'{�?`p֪�,�q�c����nb�]��ω����J�ywA�����7A/V�A$�_�<
��\��=���媍>��ڪ��VK�,rkH��X�k�/�<8Z���k�<J��^k~Գ��Efy��g02xlf����l7��r�Bs#1�@��9J���ȱB��Y�\�2���C[���<�f5� H��s���Ʉ�������T��)7�ׇ��n����1�e3$Q�t�_`��gЗ�}���/��ϰ}���%���`��	+�x��$�v)9J���X� �Mήf�ך����Υ��ɥJ�p����`b��x�X�o� �C.���|���9#�6�~��I����w�ک�3a4���%�l��L4c�\"x~Vd�WS�.�ptЭ��K���xn�Y�o9��el!o�����(��2����$�Τ�%{�W���ε�%v�QE�K�\����02a�[4%.�8�:셅g�~61:A��Z����!��~�������9��E�x_�r�V^�����-��ɇ#�֎��)�?6J�� ��K�;���?�;zё��`��	���eh�?!gf���9�T��z��d'��1�� ����x~�BQ�Zj�E�f;��s�#2�h=�_�AS�cU����Ǔ��O)+��2%U֛KՎ�7����׃�J�e�G��RXm���coA�5�X�q���I�	Qo�@�w��1�O/�|y����x�̇�+��:)����}��(<bhkTR�1���G9T��d	*5y%e숋i6���T穗R�7F���1n'������o�E��_����ʢ���%�L���F6D^Бyl$o�W���(�h�Ci��R_x�㡥/;��1{���Ђp�&,6\����������	�{�CݎƟ��ךf�{�����~���#��E�����9�C����!�������;5����m��!Y ��}$�%�[� �Z�� Ņ���9v�%���<�t��B#\M��)iR�kf
�z4G6��7>�fBPmF� z����)2=��q�w�U��u��m�P�4�V��k1�9�a-�/1�A��T��3H�!M*�׆re�IpX�Qh�;���5/.�����s	�B�&D,���
�0�>Ў6��1ƌ{(��z�!8����S�Ki�WLf���ԙ�G�{U�FQ�IFl[���(��Dv��6R>P�g�ܚ=V�r�i�6�'�G���R|C����Ap01�r\a~8�;b9a���7�����	Tadl������{��Sd/�r鬏Q��/�ju"g?c_�x0&ë��k����"8mu/kh�2���=�����!����IǮ�ԁ7�{;��b*���׭��?o�s�����ZZRV8ӥ���N��ا ��A�6� �cMJ���$ C�ܲ����З}��l�W �01Q��W��!��㫓���(l�:�@��	��Z�����u����O~�.�u_e������l��u	>���[K��32VbP�Fջ:a��eD[O�l�ϱ�	"�R��L|i`h�$A�s+b���2Hg $>1�aF�ʩB����ṸvJZ�E3N��Ԗ ц*+����3�ܞm">C;؁�L*�X�$J����Κ3���tK���V���[H��&��nf�.\YA�d�'uG�$���|W�{vڡ�EvGaz��bA�N��$/#�wL�ӫ�ĚS5m�Q@ ��:gK���o�$�i�
��?zҢ��r,uT��GMU�x�.�"9�#�V����Y8R;@ �5M��9Uz �a!E���`=�sy'��{>;��;I��|-�g�D2ߝ�o.�%�}�͎"�O��^��R�$�?*�=s6c�)k�0'}J�̦Mf�����U���Y�ދ�]K�ǈJV:�_������l�ߛ��F3C��V4q�o���Q1���Ѱ��@�P9����L`��s�Y���GC�".����
-�[�5�h����F�?������}���|�	/�$!����2�PGgW
cs(j�Jۯ�9�6��%{1?�@D��oa"k�B�NPX2Sx#i�BH߽�Zkt8�d��	�O�ǔ��.'t�\z��nw��������a������L��vlz\İ�t��s1��kq��
��1��gE�FˁBQΤ��@�-�lG'��b�����x�Ckަy0�<^��D�J�h���Cfg���H@���Q�_p�g�d1����8��?��+sE��7��@�tLA?����(x�.V�s���&��}��d�kXT�����R�;��-��h>���kZG-��~�e}�A����q�s�7�t���b�my��ZǬĭ�V}��w�7��^>޸z���&(��Ȅ��
��k�.p�-��m*����%S�l�u�#aԐ�c&`��s�_�`��.���?#A�j���n���፺[|�ؼ��k&����H���m����H޾`4}>�j�/W�-z�8qI��k�0*�C(��F���9�ʣ�Fu� �����8�����xY�kߔ�p�N�B���j]�r��a�T����ֵ��B?��vlo���g~=�AP䯁�����G����>o7ԆH�u
T�ί=�� �͜n7>�b����Tzԟ'C�{��E�J0a%K���'v����w��y��#g���lRǺ`mI��ѫU����>�����i� �6K2X�<c�������=��TE���x��H�%ս�=��U�bTT����p�3�0��ԳU������m�񽨞c]tC_n%_��(L�҉7��?a
j�~�.�O#	݋%p-�$y�]�����Q�KZ�j|L�g�����ObY��
����d�R�c�|'\P��A�'R&c7'���;�aaZ64�R��U����m��,�� ��3�����״���0����z�Ʉ�p˶-2gwcv�m�S�MMr�B��WF&h�B#"1X��U�5*����b�C���&��ߍe�g��s���ai�@�'}�&�������������1{PF�h9�Q1Z��yg�Y뚀D�/�M�@�_��|�C��DY�]�ܦ)/�P(*�Ќe�W�����Ⱥ�B�5����#�RJS��uW'̱ �����z��gҿ�>~����"l]ݪ�h���M�ڋ�4M7�fK��,6��O��b�q[���
aҡ��6�`V^��CA8vG����#Z�ԅ�1���Y�yqyG��ƹ8���iC��,�?s���J^ڌ�B\��Kd�]�xV�ܟE����4����q�O�`��`�V9�O*��
� MD�ys����E���a5��ڏ����[A!	4�<��*�'�ħ:t���8�o�>��-�r�U��.��K5�x��V�,~	{����?"�+��p�<������[�V�ao���h���P/t�NV��,�,0�B���wi����s�-�Ӟxʟ\nN���򦮰E�/R{�|үC��N�?��c/�1��/���v���f+B�$�U=���A�!��R%��s_cx�/�}	�mK
�;_�"�I�ҩ��T��z��Wr��n� ׆S�p�\�&���e�F�Y	�Q�I�M����^3��� �ԩ�8&��y�/�H>���@��L��,��1�� ��S;�5m��}����j��wm���3������s��� ��+ߎ���5`3�(<]�~hwJ� ;� �������2�#���ͼ��&�YQ�q"1z��G1:"��{�p]l6ޠ�N�Q.!B��VC�G �ng�i�_v�� �]�F��C����E��|����I���ߐ""a�����ęNvIq�aˣ�ޘ���P��ج�DG�/ه#�3zB�8b��3{dXׯ��i%8Y��o��1)�����!���'�h����;Cu��%���|�w���r��I�x�<ǚ�s�옭h�M�Xk9̱J�GU�9Y�Z��v����zQ�vI�؂���x3�"S�$��Rt$G�
�m';ܻ�)J��e�m����g���ϑ.�콍�%�ɎjB�ns������_��Ҍ�����n�ƅ�uU�]`�#s¹o�?���r��0:��X�@s0�ww9���&$�@�C�����8}E��B�޼F���W��Okk���3<��r�wJ����O�ݫ<�Kv�U�:S��^W�����c��H);�F��J��`z��pjF?��=G钰��S�=*:�3,�˪�%���d�pƻL��p��&��P�*��d��D2�z�b�6�w��P��R�U����y�n�k�G��P®[�"GlS�&��ӗ��D�CAs���Ə�V�������kDc�4C�~^�@$Z��ۙ:K�GX��Uۗ�s��9�J�� '�R*�y��U|j��!�l�q�T�����o����9E`�N�v��a�֢�F<|�{�N�G4O���]H�XZ�[�J��;��[&��R'\ ��y�t"insޚ8�Z7P�c��	X[{�Ȗ
ޮ��C�^�	&A�C�t���8����E����m؈��L�lF�0!*Q�@R|�c&�?|������M'�d�k������Ir�"�o9&"�@E�R��]0lV�u��ъ:�c_���ԇ=�+���s�a8�0K8(�Wyt��@�筄,|gs�RV�u8��s�q�u�Ù�gJ��*�@v��g�4��g�G�X�*���nj�fJ�u�B����-���M&�-z&P�)�Z�	���q�xov �Y���C��@�Bzi��+H�RL�E�I�Y/�������M=�M��?-�{c2@�2ދ8��mU�D�qʣx�4�?>�ZJ~�)�.e��=��Qq$pJ��N]���P��d�cT����w]Q�j9�dp_5)Vr��*�>i�b�ޕIL�=��}�HG�2�U��$��v���8r�Ț�O�$�\:�#�*�S,bv�óxPN>_���֥B'f׮�(�_���%}w�؊@.�
��9u�|2V����\��Ų�����YM�-9n0��'�ϫ�̖��*�ˊ�~`
U�W���kGu�����V&�(ɫ)������"M����dX�l�˼��W��U
���~�f��� ���2�;�������5��ɀ��,(]�M̀;��h����_ӯ��ȍ#�&�(����g���t>J�zc���3��:�(���l�bQC<��9�	�V��c~7dV�/=P��e��J��$=�F�b:�K�#��d~���|�~��zd���x��ź��;X����8��v�㞕�K����m�Av�^��C/��UU� �<����A"&�Գ��cR�����$C;��o���X,`8Gp4 {����(5�߶�����'GJ`��,F��]3�<�Ǧ����ᙳh ѧ�7?C\$���Łx�Mj��a*��!�J�����Ս���ߒ=���:��	�'~���˓4	�5eV�b&������ƭrmt)>ݪC��l=��|,�]a���W�n��᥿ ����k6�f ��zQ�fC
��{�/�ã4aS|~
�w�G�>q�+�R����~�n-؜�a�ħh�b�у32����Lr�k�\�M^�xI:t����5�*5�M��~�Gt�i�Ng��p��
p�L�v���U��H���G�(R��WA����r�A�`���]=Ԯ&oXP����}U�kq7��D�l�X�d��A$o|�^�	�	�߾M�ܿ<s�j5ŘE�o2B3�N�.M#�pQBq����<��x�����vZ(?���R��1�W�Ko��Hkǭ���-�A���F���:��(dtX�S\r�A$�d�p"��+�R[�*���٦��ԯ����^�i,F� fo�=��_pI-����i���q�,�#)_�_����/){R���gk�h�9T�,!ȧn9���/F����;/����ؿz�%��0pÞf1�LHP.���r���儗,;,*Q��.�qc�������0jyHp�Ox��)p��0�SP-vA�3����៚����l��)�N����l�|p�@��jE3��X�-���r��T�|�Q��: ��V?�v�i��W�c��/TJr~r7��l�r��-�h�a_{��n�~n6\.�<�!��
�ϿJb��^�13�o&�r�\�ET����bU� (&,=$/�8��զCcj���ej&x�gdc��q07Z��!�D���r)1��N�V�m�����*�씬Y�X���6��������o�`�a'��&�ӅMΎ�<T�YB\��-i�5z�6p:-�/��������-Ny�$�����8�L�S�vXI�c1��1.�?�J�G[&�K�~h���E����;5-Fj��6�I"-z`i�%rr�~j�~dug�k(k?@}����ܗ'9�գSV���k ������T�"��e����Er4�c�Z����\��#D b��g)�	���s���VNm�qe?RY��Aq^ /M�de��������~5�JI��x1�ݴ�F������	���<�J�u�)��*���3(�]�������˿�F	b�9����Po��s��u6��������?GG��ňR�ܲ�3?S�i�.F�,8��Q+yՍ�bG�V}������l��u!
<� ���p�m���j�Oi"�R�4����!�<k�R�����lպ.g⮺v��_9z#x⏼d��?���T��d(��X�m@����t��_������1�t_G�z	�<��O�pl'@<���Xx����&���;*G7a��j�Roi�*Q/Hi�v�[�?=
2@)����X �H9�j4!I癘�$'��6��K{������7B6n�L��«fK��4�~D��-�%Wi+�Sa��ȉo���u|�������TU�8۪|ϓ��,X�V}��+��K�:�$wiYHHkn�e�T��m6>��2!,� ٯ��?ރ��2�w�lGDc���~ڃnx��Y��KI,�?F
���.��A1�����o�#�����(9В�kd������|<_��el]|j�����yv�'^���h7J	�{����`��`#���vvU����F�zE_F-�Q�\TZ�v��QQ<M��)�7 @٭t�
6��8��L1�MKm��l���Zn��S�uJ���YD�z�ϲ�,B<3ȧt�Q�3>�=,/�r;k�-}��f�f� �#��#*)���v!�2�sc/�9:&.ʐ�Fr#Kp,�:��(2'5���\?�Ъ�jIU�.z�ո�\|(N�涤{ �U�$]H��}�R#�&��A~\��Ҥ_�1��>j1�q���6��_�d��l�XJ롅^ސIG���}���ה+}�,��=��I����
h��^�課��6j�OŦ��E�,�F'�Tk��j.������H]��A��yNw�YEJ���@V��ސ| ��!ku:�@em�J{Q�M:6k(?3�@z��T^ޡڳ]�<D��8��eY�}!
1.�\e����X�h�A^�	.��Q�|΂����W�@&xƏQaM�Z�h��P��65�K3!oY�S��<��9�j[�I�	��AԅҔ����YzG�N�����/.w	��:��<A��/\be7�V�N��ů6��/�
�Ȕ@�ړ�bS��TL�Ի�ު��j�����w1�,KY:���䕑49S�ZK�����ډ
,�(��Sg�|�H=�°�ˢ�I�Tr�Q��Ek0�B+��h(N��j!z!�r�9i�ת�i�G'ַ �:/�49���9H�@3=�6'����.��"�����-`�;21�o`H��T<>��4[y�hN�t6�����Xߛ���s�͋������7�躊p5ҿ�46�ҋ��$�O�����B�pR��?��� ���Ϛ"��2��k�)�R'c���W������r�X�,q	�+h�'�\�����UHq(f\���7R��g��"7�u��{6UŬQ�N�`73���f�r��T���g�,���Bh���h���r���f$CE���R8C�B��v�<�e�⤃�\;�4�6|u� @�C@uc7�0;D́!��˗��᪍\��g䲎t�`��{�L���z�󴸰�~�Y���bj?0��ݩ�hM�~Z����w;�$��.+ ��_1��;�%�@Y���dVf��	�I��4�b��kr�% ucԾ�����gޤH�������5!�ᷛ��G���vO��3Ƣ���)DTI�؄E����,e����O �y��A���Y��*��I6��4 �z��t��r��6��� �֝\tHF��:԰g,xk�s�r�=�s��SICSNߥ�����,>���`�)�Ӣ++ť�g��]��@z�<5��X�4�4l���r-��)\8�F��o쒎��rW�	�(�Y4��j���S��ԭ���γ vᬌU�@�_&_��Z�
7�� Z�]qV���`�M�8���T��_]˛��js2��x�b�8��#�M�%i�Y��=!���B
��ڨ�� ��I[lpFnz!�	]���i�g��gr�M�R�w�O�'��"`qy�P7����D~<3!A"�\jn�? ��b���޾!� �c׬�\�����"���p��QH_F���y��V���@��5$�f�y,lx^�Tn��D&O�J�ůZ�(�������:E�A�jH�Nd6tK���:�LZr	�W|<��a�M�����ׁ�IǺ<�8�wP/�|�R�	"��  Y�7���Gn�S�Pa�Y�aؚ���:��y_���.��<�&bm�B\�vH��_��ܐ�er�����O���ܥ�s}N���c�4<��Bn�n<^��m�sБz����a��kl�Fn�E�����`A��!�1��eX��|��|�G�Ц�9(Tg���T(f�X����wzQ6L�	ӊ��ľ+G1��[��%����1����K��m��s�h���`��[��~�6���bGi�C0m�%��í���ɴ�^ړ0j"�-ùG\@#r����CO�_!s	�%Ca5g���R��5���0�t��?&���0�FK;�ڜ�D����_C/���S�ݗU�l)���7z����Wl��LcAvY9�a��+�m|)ƒFgs��7ߏj3[ v���@���3 ����X���~�(3����?�wG����.�2,�χ���'�[8I��)n��s\\S��im�uA�K\�H����Zve�n�����R$2ʁ�BdF�=�'�˱5?0O��.D�3���9�{�gP�;U'>L��LՈ��3$ee&��Ap@�M1�Q��*�6�e��@����X�n��p�X����� �p�&xU�7習�h���Z�dU��9+���i�䳂3b�_��lût�j�t@IP����-:�E}��!���$���,�sVn��#1��-��a٥�R����~=!LR�O_�(#/o=4�M�WRL�Jw�|�)���{'��.��I2�9�"�4�?�쟃/��˨I�b����+�¢0�AY��h�+��8I�5�j�Q�dVp��]W�3�Z����.��f������1�l>ze���\#���׈�����˃z�..�ǃ3���'��Χ�Oj|7�釦�`�v�=va"A����Ӵ�f}�2}<�,�W�����IWs��'�Z����yR���VHԂ_�GG$:��?�*zu�U�d<)Y��l'�7B��q�S�|�K�DH�'^�T	�)8\�������ؔ��r��J��8!g��u	��.i3�sx�ض��(���b1�p� �"�q��'��Ex�`��\7R�>�=��(_x[�j�o�ҁ��������]�Ѩ�-H���Ϝ-�ܓӗ5���OE���znW�ӑ_�(4�s\�z�d	�bM�y1p��[��H"N��&�'�,a ��O�{�{�"��g��j~}���W�Dl{�ɏ1-b�V{
x�q��T��Ǩ��"���X��d4��U��#&8pl�Dt����Qֲ�Hg�J�V
�9>�՚X�)�!J��!s�iP�����Ɏ��J����/u#�*x�{��$����v��+�$�2W�ԋ韟�v�%{��C
�8�?^�&֡�呃��F����n/����\�F�p�@�n:�&�xY�Mܘ$���}�:OC(f��2&.Q�a���v�-d�޵s��<�������o%�8�鰛ㅝ�aLk��A�)�!ZD��M9�4�G����CBOB�tNF�(J�>HXj Yͼ{+��W�����dM�F���?�UeK��!0\�21�E��`�
u��sc#]�,�����KBF��*�ʠ��ѷ��3�f[?��c�(���+��{u��v*�F��f�m���<cX@�5�z�e�X��r��,?��/�R��3#q.\� ŻD�# h�v�֨j�Kq�p��4�<���~a�)te�ٽ�Ի̛�)X��H���S:0;�4jB��kO�£��]�}� ��v�q��_o?�x����jUP�ՠ&�q�'��|��(JCU�Q��_P�ɢ��;Y��q��� �|�`{{5��tcӾ~���B2 v�3�~�ThM3�M��F`фHx����7 Mt��{K������[������Q陝���~���	����a�n˟�� ��h�T;��J�"�g��:�y��-Z��,���v 	E�����&�Cn��Q���F$̒�����ZE d�M�넹����+�29�I���"Ժ��/����іoQ�{KQ�}�U���
Y�biDC�B�/����eXj�e�vh�G0��y���)��A.�S�W-�ω��\���/���w�S}���F����ے�+ǅ���k�2�y��]��W+*�'�H9N�ɠ/����&�2�<�->���}'��F1ǟ������H��3���n{�c�����)�n�C�p7M~B�l�VUY�f��1[R�Lݚg�J3�2ָ�LN1Ȯ��U��&WfY��noϾ&��Ϣ(%����n�O���� e9^�Hn��h�~�ܝ��y���W���9�g&A	�N��4ͤ~�̹IDA��H��{c��8���I!/C���0THGP*����^��BX+T�O��ƺ�r�,@%%��#�o?uTfZ B�´%�A�Ɋ��h3�05����1@�}:�������S\.�2�"�4�`�?Ϳp�����
�9�vCx!��|��i�ñf�`�����!Ў�X�*u�+D�[�^��;�^s��#�0��'�f/�� 8��~��<�,22۹��Ȫ.��ظ�3���Q��uj�0�V�臗�A�g�縃/��ѫ�9Q'7�l%�M�bg��u��2���*�n(V��X���R��;�@�kty����j���t�O�1X����
 ����0
�n	�;��־t�|{�����q�k-ýk1(Է����T3�h��I�'#���M�\�)(@"�8z?q�[�p|�<ʋ^����0$ij[B���q�T�XR͐��x�4��rJ��9�+?�Z.-Mũ�ɛ���A��L���_�̠��."DL�蒳t��ɫ���0@0	/��{��UƲ+���޲���a��o:�?��&���oH^j)��"��<Wl�v�%b��}Jd��,=�'��x\�T�����$q}͎9�K� |�ӵwC_ԇ�G���lf<j���x�l���+b���! kW���2*;Q1��	��.��ٽ���_���3�Ƹ���T�^�v�&;�:۸<^�rncZ�ȸ�L�������������D�zrH��Wɢ_y�ZՏ���=C��c�֯"�n�R^���7���}.d�f�Ɩ͹��wV�H�̴�V�X�0�HJ��NF3��C���g�C�U�
w����K��m�
�Nlr@[ݏjځ�a�X��Ĕ!8e*e�v��>��/'�`������|vʚ���+�|�,�.ؖ��$Ыܻ��������D�;�=��p<��-����Ǽ���7�n�J�N/�c���8F��<�}6�`��rfC�1!�!|��\9�ۧ����������=�!q���!MKE�5_9��EW��� �G�0Vɬ谀�
q�$J���c�.Yǹ���������6��&qt�fʨ_�HR8s���Sp'�{8�K���x��l�`,���Q�o�T����Eڀ��@.Q0f�ɡ�!��M�`\�����W
E%
Ԃ�A�h	��M��c��4]�{A�N}Û�%8��]Oj�����~Ğ�U*gНc�oOF�D�J��v��:�y���k١X�B�t�5������Y��0^Z"��>��';��@�m����c�T:�A������#x�es�>�[�x �8p��"S�7G�:
Ly���r�R����tP?x~�ھ`����Ѩ�ɾ��G�p@�5<�������$�Dz4��ўc�DHy�,�����׃B2L��ica���~y���p@޺4PR8�b��x��Y�eV=���lo,uK������9�l��6�P��9tJ��3������aq���#n4��m<�<(p���GV��b���p��B�IcG��i�v���Sr:7��r��rd�隇zED���,��t�����Ƶ".� � *�ё�O��ǐcT�5$���VJt�ɱ�	M�7�ӹ
4�~72�H�?TPo��&�e׺k܀� ���!���!�`��w)gI��^8%���za7W�}����� �Qk6����,l99G�&�(~yH<=D�@-
WR�G%�\-��H+k��!�]kg�d�N�n�^B^�b�Y�
��U-�}� ��#/|�X>���8.,�7��^�+ٲU:�f���]�v)Hg�5�pf[�S�x��h��7N�nժjp�G��ޑ�+�c6 ��e�p�H�ӝw����?'��� 7>ll�w h���f�u���)wՀՐ�����z�V���.��o��a�t�z�~�#Е+����U.�K�� ��S�/D�P�bKg�D�-g��Q�3�]O��p���)�1�8ldQY]cu��?�=[hy�O��R���
{&��\�"����/G'��\m�n�5�+�U���M��'�'��1a,m��H�}��m�U���z�I�O��+.�N١��b�_ͩf���1h'6=a8�8����������l������UW�%r�K����T�>�.�OV�C���o�K+�&#
FymU���T�Io���Չ��Q�:(��7���5�n��ih,< (�`�+` �:�A~��80�p�2�%�k�������9p���	W��#X�F@�z}��@V�V�E<��Ԑ���r�Vt�J;2y�~����#�>[e�XH�Q��m��[`:�`�P�_cr�8���M��Xah� �N�^����[�7u�V�׎���Q�8%���f��c9��=�{Ʀ�X�y��p�K@��UPm�r�U�ƫ�����=uΔx�"��o2��#�{�MNf�D��C!�&�Br��%r�0N�դ�aCu3�%��ePV�m�T�3>��}-���w\[����)=/�_�f��H���~ �*���i�}m]���/_���8{H��M�R��*~b����xT�TJl*u���3�UȦ�%�b�C�����+~��2p)Z��a�Ʉ��Xn���c4fd:����$>�}��r�"\Pr}D/�)O�҇966��$���o�k|c�-)]+}�6���C�:0��'�*�|+�O��<�������C�c?��9g{M=D��Jp�@ �4X�[�Հ��*��'P��3wdQ�Օy[:,H�g��~ܖ�YW�̬�[]r�7崒b���Ѭ'�y���2l��[���I�߁j��A(<�#y�S�蜳���ǿJj2��K._��%�C��z����ا˱~�l������'�:��y"Vj�<޳b�&�jWL ��+?�@hP5$,?nғ���7$K��N� $d�KĈ(d_�zݹ���� ;�����s�5�j:@	I��spZ���p�,%�Q��ڄ����z���$ׂ��E��1Ϗ��m����G^T>�����­Xs8�ȝm�l	1�^G���1�Y�����%�- �Dt�X�f��u��b�	_�C��ե���C��!��ֻ�ke��;_��F��\^�[�/���e���ʅ���S�����
��̣y����V�H՗s`��`�7���Y ��B�R�O�lj��������@z�S��$�#���F\��� B������EwLg���CP�{���T�E����_��">�:�n�;VT́�q��R�C,����X���#`��Kغm�)K�����M�<��~�R�2l�wJ��l����f;���t���pg-E�5�C��w߫�{~!as[b!���0ޓ�^�].6���d�*���Nڍ�l�w4$A�
�N�/8�u�-"����aUD^]�������e��	G8����a�4�)Ť��B<����	k��9���^��(A�P�6������\|��+^9Z�%��D�\L��+�*w�b(;<��������ʃv�yĴ����E�N(!h�f}$E��3�Ed��[A�����Q�4�r��$pu=������gh2}�]��,_t}��9x����w�c;�g�B�,�q�/?	�h�`��{t�@	�Q���x���mSB�:�Î���uj��1-8������v(@���O��Jײ�3OL`Y���1O�J/4}� ��嗢}JI`ц���|��K�Ӡ�����À��L2e�1�����:W"zf��R�\Ƞ���NSu��Y尢�mY�~Ǭ�K��w�Eܬ�:����|y�=��8I�ڧ)w�V�+Ň~a�LGEf�cg-]���m#�#hdY�]|��5�"��lPFj�fAmB�xy�ް��{�|������+��/���<�ظؕ�������}|�'ImQ��(���x�8�j@���I�S�����w��i��,�nM�@g�vo\���.��!�_敢:�I ��4_(�ϛBRC�W�ק��q���Dp��<˒��{��ǡj��Dlm?���� �e��q��Gg��ǿ����y��D@ϕ\��C����=�D����,�`�M�P��W�q\'�	c�~��ð�Y򔝽{��&<Y��,˓�J����&�Ex�}�u��f�'��0����w�@֕K����Rk��Pg����Ԟ�4�iZ�9�$��(?�H]��?-�k_ՍD^k=�R3�0H �Ǟ]��Y�}K����c� }�����U��(-���͊(�U��e$���
T�g`q]��(�p�I!���� �W	ˡ�( ���Q��$�?��~� q�{���t��) �'=����� ��Lȋs.� ������u��n�]�gO�8.$�4����D�6q��fR�E���U�}�<�-���&7��B�jSi$RN:��m�]:��SI�Y�>^�E���zd�J�n���<�j��3��GKbt������s2Л�"2�퍫o�ёV*�vd��(�ç�8�GF�☾�0�P��� �������X�&��$X䆀#l'f���;�� eo"5Eq�.~XXf�(�M����M��s�M��95�%�����{�DC�단�fpݸB!�7Ub:4����N�~�ޗR��ŝc������q���(+ ��a�	-r&_jbtT3��)�1T}��2�<Q�L���[]czѷ�#W
G��|M\?r�bF�L�_T��n�DC�E��J��!�k�:�Rp�T�O�cӢż�g������0�3�N��-�iyӭ�v�VN߆�m�H6�����X,�]<��LV����،��>U�3p9�y��f�b��q}�yLVSѓI>�&@�7��wX�5d�1���<�:�!/�z(|XSX&���j�W"�@K�H�#ȥ��W��p̧AF���!�ƀ�s�v�el0AV�T�u�9"��v/c�CHv�!W7�ô.�ʜ�<޴�(�/��X(�]�^U���&�*��F��/���������O'��5jQ��/�k��+���kw�!'x81�>�c��KPЏ�KgTH<�h/��3�u��/p��N'�v&O]�@S���/�M�-?�?�Ҕ��-�6�x��gM3'>"��`�^���._�`��:`����5���w��\�`z�¬��y8��K� ��z��7�Z��D� ��E��9o�����q(%��-G/I�4g"�n�y��$��w�)*��r ��a�i	���P{��/��<��w�췈�Q���J��E��j.�8�"�pF,Z-� �L6�#�T;3�ڊ-a]gyVF�8�%ә�Cr
�
�O� �:7���T}NH�΂��n�'�f�V����^a�� j�O[�S�ˠ�\��kA#��z�I��3�s5���*�P�����5�+l�f�a-���[Ձ��(Z7��G����	D�����$���4�eG���(]/X�D���Ap�^V@�C1�W��AF��c��z.�PC�B�Vr��J��;�-+|��8f�>��e���]��� P����ʾ��\ eF;���۷��IS6F�H�]�����ٸ~
�a�����-F�_x[�G��j�^��`��<�	i>��\N��_1��_�D�-k��{�VR0|V6X��@ij$����V��)w`����~4�U̘��zr��\
��:�r�M3�[�M��2�26����}�'���%��4It��3�<{M$��tV	#<���&���6뼈r��&�'����\�:�������v~�R�,]�9��G����+�n�K��4	\�Yju?&�`����r(M�,��L�t���`5F2����VE���jW�zq��0�O��([γګ� }��j����ѻX:�\�}'f�+�P�"�a%ۗ�81�\6��/�j��Sk(�|��y�������[l��ӄC<[���P�]�.�(��[
4 c�MI�-�Hov�}F]*
ƉKXȹ&�H��C�����S)1
�>��/S�MF��� l���0��T,S|�ďݎ�nI*�,n�q; ܔQ��yJ^t`��h��b!0�x��Q��x>2�T2��]�T��W~En4�����A"��t��*��?�����v$K�n�����.�<01rkS���ۃ�1ê}��L1��v�GX�T��Dm�	��~x��(�Aeo����|tVΒ㮶%��=X�Dc������\�D��R{
�N�O#+au��]�K:=���JMF0���6�U�|JaH�C��d��E��fn筤Y��'j��A�)IՔ��Ï�8�!�J�gZ5�骥[�r��2���L�5���-��B�ƛ 
ݳJ�W`��QBN���3O�U�) L_u��1�-j�`��{BUȰ�f�EH��a�סa8DXpn<&kD��5�����˻�&q=�cT�M��$��"�`��F^{8�z���u2�F�?�	Vy�
1s+_?y�g���k�q�[@�L](�6�M�J���4����FU�=a�>(G��<K�(�)#����[�8g�j��W���{yֹh���rc@��;�ޤtᗛl8x�N�O{ܵн��qnú���K'�"3o���_!G�:�<��K�鵘T�4ռ^;��>�@p�*~�)�%�r�j�C|��O["j���X����!����m���z�u�.�^GXL��U^�@f�c����(�]{�-USʁ�qܖ.����LT2�{�9�[髽2`8g�i#�e!��*����ɵ��Zo'0�m��B�7�3&#_���MN4U��k��\t�[4�|CN�-[�������G!�[�Q[
�N��e~���	_]�[�^�����Hn��{&m������96�!ɖД݋��]��n���汎u��U�bPƘ�&�3�g?efH���*���Y��u�PY�~r�t�i^��u��{�#�d�ec(.p~@S��I�9_m�J�����b�v�;tM�1�~�'����./�9�*B�Q�Ģ����G"���75�e��&�o�g�uTJB�I�x�۫v���:[��}��~4x���*6?�o{�,X���Է���V�h��ۉ}!�b�������Qt{���Çe��e�{���8Xy���mCXLC[yG�0�4���W��y�i��n ]K� od�;-e3_I�{��M�|�_�.u*%1$L7��e^�e�I.��i��Js$�-��B���Q^�������/=+"ݢ>�ɴz��`�''�_�;�Z�]�oIM��f��,���s��h�o=�G�Lb81D�k����N㟯��N��L�r���Z�����ž���/f �D���Uhe��l�[�1j@m�C%��d�_l��4��Ʉ�8yl�����FA)�?��]�e�H�rY�j�{r�?�����Q�Y����v@Tl4: L�j"�_{*�*���Q����v�s2�x`p�Z(���A=(��)�m��:���NtZ{xm }�X����1V�jPԠz�q���R�b�|��@��`��7K_C#nVm�Q��v5�-��ۍ�ĺ��Z)qa�zn��\-�����C' �Qx�\���*!�]��CZ�>np��w�A���t�F�5����w����V.�&��׵1�ժ��e��d���'�9$�Pp�1�-���w$�*���C���͊�[�9j_��5�'!ZmB��Gd8�E�8\��(z�[ه��ҡ]Q�rq�D�m�����~,���4kf��1%[o�˞C%������ɠ*�?���9�IQB�"*����Q�8�D�	 ?���H)E?X�KE��\��YŬ*�?�Caq�N�ʈ���ry��Rjj���i���+(K���r^~$K`!�.?�t���,�,�s���fÚ.ǈAqvВ��^\]2Z*��#ba׹JT���U~�]E2J�h��l�����-�Y'�����[�ki�+�M�/��p��WE�)�z=$4���+��\׽V@qJL~�6%�3���S�����έ����v��B�[+�HOKBS��jQ�`��	��&��s?M��(t�N����~�L�P��BeGb���U���Z�2�R��P`)C�ΫԺ��ua�����֧�D)�q�!5�բ���'�F~堣?�Jw!��ůs0��x�{KG+�Rl��i:��nl��h�%��+�3��M^(Ý��kC�æp[�5���@7��5O�� ��p��G
pV�:x�I����[P��R�Ѓ��2���1�S܇�Ar���đ�,kx�q᧎A'�IL�&�:6[5ɻ �X�c����!�n&���h�C��@�v����Y��' �[��£r���;(T7hfLq!��^�k�l�SO@dvo����,u�d[h�{6U���꡷�{7�����5��&h�z���u����B;`c����<�G��eE�?J�Ł^$�VusW^s��P~<�N���h�{���n$�|V[�0���i�ҶFqRp	�	` 5�K�,O��U��q�HTl��;	w|��<GFTOm��1�$���ѻ�~�~]i"�#oa٤s�g�����P����Q`��T��(RDX�T4�m^	9�?�k$2 =���֟�zc2�u�F�"B�`.�e� �,�9x*1���}�@h��	��	�=��G��2;��O��[G�v��A�S��[6�BZ�V��F�=���7�+� V��Z9wEt����熋K��;5[� �]�p�����&\�ϫ�h:��֧���W#�-L���Pʴ���&�M�N�"U��8kK$ e(�;+�T�qŅ8���x_�hT�x~��~B�c�n�*��F5���]q�h�qfX��o�A������&@j4����˳��.�g�ЊP���|3����Ȍ����ŧ �e�'9��~H��,F��P|ԸG�̭X�F!9,_�\C�i��!	��E���I硳⋋�D�Tݐ˂����kF2���
[U��ѡe2@��h̀,����==�-X��d�$?4��|lu~y$� j���^0���ȩR��[K�����@+��<�ꍝ&Nxg��=K{��U�4�\���WEؔ������)���XQ�W������G��l�[>4����/�$d"�;Yp{Z�5���?�����6�;��g쪌o���D�B�j�d�ʝ�P����ď�v:a�c��jeX1���l3H��g�<�����o��?��ڢm���8�#���90���ȁ2��c�D��T���o��%,�kW�����i;�y���	{"xf�����} a��N;ި��ɟac����[>7��́*�e��E�|���L'�G�U�چ�	laρ	f����4��&��G���f�K&a@�z�S�x%[�3öx ���RK`h�K|����J����?�-���sa��L��vG�6E&ҹ�i�m�M���z`�z����Z�<�Q����z1���k%��dpdӓJ���j3,�AVxS�aMF#��Q��:3��� Ү]2�����A�Lzh�~��5�w}����,޷=���s.���e�t���X�j{)����K�e̽�cx!�<�^R���>�]gw@'H���u 1x>Bcr<[T�����Wޫ��I�1<�������-�C`���<?��]��/d�d���7�v�}����J'I\���JJ���S��TL#�FR�wQO�Ĥ��h�W
���g=}����������?p�@w�.mZ'B8b��l250�5��(��K!R�Y��l.�L&���A^N�"�D3��K'����d����~��M��q�jLmY �6�?����#ށs&��˹����٧��j��y/xK��45����'w ����ŊN-�r��<�~�:ګ7r	��U��'�ua��a��668���D�ȸ`ƂiCd�s`%�{k�!d��Z9/�e���E\1ƢK]�r��#��eu��7���Jq��DD�ʦ/�v!^D�T���v*�Y�C	~G�?Ev�8m�u�,�u�,��A)��J���y��e՜��ݺ�[Ԗ�A���?�T��5Ӯu�FË�/
�lU�g{�UDV�����KtC\Px�r	?��r���͎ײ!\��A�Y�Ȳ�ӱ8�n���Y"u����{���x� ���V����'9�y�lf����s��*o��@��{˒n �g�U%����Z�,�P�Q�g2��8��'LS���VO�
WזM��j���;ȭ�b��A��Tq; 32Բh�fwX�;�b�m���'#�FS�%|Uݯe���{؅��m�W	�C����߆��yb�a_V�<`���F�'�*�+zʍ^pJs���w��ݒ�;'���J+��U�\��[���9#Z�+h#�/L#�]���@$�p���r�|�e�.�~pP���[nI����/�_�#��{MXv�{u�!U�d�u��`lAUnL��7�][jx*�|�x��i���ۄp�z�����ɠ��	��ؙ4��G�ԙ��OU��ҽ_��F`q��o|��� ��_�FKg{�;�'C�Y�Fpv�}J /�q%G��E�皟�4X�y/���u�mX�N5��v�R!�I���� ս]�FO��p����Z���c�K�p�<2y
��#�Z8ꮉՎCE)0RV�/ѿ��*:Ȟ�jH����X�i.IKu0�Bjj6�rc���1zU+吀��id4p�	�_;樂�O�?h��κY@'�g��i�>�cãm��ZY�a�n>+�0NƓ�ݫ�1�;��v5dr� �0�~lu��1F��haY^Np��-���3��2�P)
bj1!�s�� ������K�'&�ZwH����.�%�ƥ_+����(�L�o�gٶN�*���ah�"Z+�u�?:��a��b�#t���C�c<G�j�ɶobF��<�����Ї;��l��KXZ�=2.�v��������y!���w�����Ն��Ξ96mA�N�4I8&���m[Q(Rͬ����?� TR�r�1���E�(�?{�_��4�{���@��"(�Z��ϯ�����[�^.���,��D�RWfc˓9�ytzO��N������!0]�F�ݜ��<�q>0�_�0��Virw���4��	ۿ�I�(�i��l��59t%-<�^�=�k��-.<[W�(M��IP]o��'5�:�J�aD��nqFl��MZ�ϟ@#a�^��%
���8�D3���C�dz�� �
�XF    r_�6          P  �    �    �   X �   � �
   x
 �   ( �    �    r_�6      	    �  �   �  �   �  �     �   H �   p �   � �   � �	   � �    r_�6           �    0 4              r_�6           �   81 4              r_�6             p2 4              r_�6           8  �3 4              r_�6           `  �4 4              r_�6           �  6 4              r_�6           �  P7 4              r_�6           �  �8 4              r_�6              �9 4              r_�6       0 �x �H �� �X �� �p �� �� � �� �@ �� �h �� �� �� �� �� �� �� � �    r_�6           �  �: �              r_�6           �  �< �              r_�6           �  �> �              r_�6             �@ �              r_�6           0  PB �              r_�6           X   D �              r_�6           �  �E �              r_�6           �  �G �              r_�6           �  �I �              r_�6           �  `K �              r_�6              0M �            B B A B O R T          B B A L L      B B C A N C E L        B B C L O S E          B B H E L P    B B I G N O R E        B B N O        B B O K        B B R E T R Y          B B Y E S      P R E V I E W G L Y P H           r_�6          0 �    r_�6         H  p�  �%              r_�6       � �p �    r_�6           �  N R            D L G T E M P L A T E             r_�6       �  � ��  � ��  � ��   ��  0 ��  X ��  � ��  � ��  � ��  � ��    ��  H ��  p ��  � ��  � ��  � ��  	 ��  8	 ��  `	 ��  �	 ��  �	 ��  �	 ��   
 ��  (
 �   P
 �    r_�6           �  pN $              r_�6           �  �P �              r_�6           �  pR ,               r_�6              �R @              r_�6           H  �T                r_�6           p  �X 8              r_�6           �  ] x              r_�6           �  �` �              r_�6           �  Hd �              r_�6             g H              r_�6           8  Pj �              r_�6           `  Hn L              r_�6           �  �r �               r_�6           �  Xs               r_�6           �  `t @              r_�6            	  �v �              r_�6           (	  �z �              r_�6           P	  8~ |              r_�6           x	  �� �              r_�6           �	  h� P              r_�6           �	  �� �               r_�6           �	  �� �              r_�6           
  �� 4              r_�6           @
  �� ,              r_�6           h
  �               r_�6       � ��
 � � �( �@ �@ �h �X �� �p �� �� �� �� � �� �0 �� �X �� �� �� �� � �� �    r_�6             �                r_�6           0  � �              r_�6           X  ؚ �              r_�6           �  �� �|             r_�6           �  p' D             r_�6           �  �k ��             r_�6           �  PX {�              r_�6              �� �)              r_�6           H  � ��              r_�6           p   � �|             r_�6           �   I m�             r_�6           �  pA '*              r_�6           �  �k ��          D V C L A L    P A C K A G E I N F O          T F A L E R T A       	 T F K V I N _ K X      T F T _ B _ B          T F T _ I T A         	 T F T _ M O E D A      T F _ 0 1      T F _ C E A R A        T F _ K N C X          T F _ K V E R M        T F _ O R K T          T F _ S A F R A           r_�6      � �� �  �� ��  � ��  � ��    ��  H ��  p ��  � ��  � �    r_�6           �  h-                 r_�6           �  �-                 r_�6           �  �-                 r_�6             �-                 r_�6           8  �-                 r_�6           `  �-                 r_�6           �  �-                 r_�6           �  .                 r_�6           �  (.             
 R X _ D R A G C U R   
 R X _ H A N D C U R       r_�6       X �0 �    r_�6         H  �              M A I N I C O N       (   0   `                                                                                                                                                                                                                                                                                #   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   #                                                  #   k   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   k   #                                            �__��]]��\\��[[��ZZ��YY��XX��VV��TT��TT��SS��QQ��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��VV��VV��VV��VV�   �   /                                            �aa����������������������������������������������������������������������������������������������������������������������������������Ψ��VV�   �   /    S,_6Jk?urD�n@�f<�^5�X0�O+uS0R�VN������Ѫ��֯��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ͩ��XW�   �   /    �QnՋ&��(��(��(�̅)��,��o)��X"�h;�nD4���}�֮���ǟ��ӫ��ծ��Ԯ��Ԯ��Ԯ��֯��֯��װ��װ��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��ر��Ω��ZX�   �   /�m(5�'���&�ъ#��b��RV�t&:�v)M�z.}�1��z1��q?��gM��uS���m�֮��⻕�໔�ߺ��Ổ�ὖ����ȡ��Χ��ԭ��ְ��ٲ��ز��ز��ز��ٲ��ٲ��ز��ز��ٲ��ز��ز��ز��ز��ز��ز��ٲ��ٲ��ز��ͪ��[Z�   �   /ؐ+���'�Ҍ$�lA�L,1                        귏�ґF��l;�uS6��cD��qQ��oO��mN��oO��uR��~\���j���y�ү�����Щ��ְ��ײ��ٳ��ٳ��ٳ��ٴ��ٳ��ٳ��ٴ��ٳ��ٳ��ٴ��ٳ��ٳ��ٳ��ٳ��ٳ��Ϋ��]\�   �   /�(���'��g�=�M,	            R(O(-L-W��~��oI�Ό<��5��r0���8�ƌ=�ÎB���C���E��v@��c;�zZ;��cE���c�ǥ��㿚��Ы��ر��ڵ��ٵ��ٵ��ڵ��ٵ��ٵ��ڵ��ڴ��ٵ��ڵ��ڴ��ڵ��ڵ��ٵ��ͭ��_]�   �   /�%���&��c!�9�P-        S-N+Ee:��Z#�΄4��:���A���M���O���Q���X���b���p���}�����ߐ���}���U�}\5�w[>���d�Ю���˦��׳��ڶ��۶��ڶ��ڶ��۶��ڶ��۶��۶��ڶ��۶��ڶ��ڶ��ڶ��ͭ��a_�   �   /�$���'��l#�;�V0"    V,O-_�d&�ڎ5��>���?���>���<���=��<���<���@���G���Q���\���o������������ؘ���c�oR1��jN�¢��ɤ��ص��ڷ��۷��۸��۸��۷��۷��۸��۷��۷��۷��۷��ܷ��ͯ��ca�   �   /�'���)�(�E&�M+_U6+`8tɃ1��<���?��;��9��8��7��6��6��6��6��7��:���B���Q���b���w�������������ň�{^5�~aF���{��Ǣ��׵��ܸ��ܹ��ܹ��ݹ��ܹ��ܹ��ݹ��ܹ��ݹ��ݹ��ܺ��̯��ec�   �   /ۗ+���*�ݞ1�Y5�C#�f?���5���@���=��9��7��5��2��2��2��2��2��2��2��3��4��9���E���V���l�����������������h<�z_D���~��ʩ��۸��ݻ��ݻ��ݻ��ݻ��ݻ��ݻ��ݻ��ݻ��ݻ��ݻ��̱��ge�   �   /ˍ2���*���:��\�?"�֒,���<���:��7��5��2��0��.��/��/��1��1��1��1��1��2��3��7���>���N���g������������ݞ��g?��hL�ί���Բ��޼��޽��޽��޽��޽��޽��޽��޽��޽��޽��̱��ig�   �   /��1o�,���9�ȏ/��v!���3��7��6��4��0��/��.��,��-��.��.�އ-�ׁ*��~*�׀+�߉-��0��2��5��<���I���e������������Ċ�mN0���d��â��ۻ��߿��߿��߿��߾��߿��߾��޿��޿��޿��̲��kh�   �   /�w*�0���5���?���:���4��6��3��0��-��,��*��+��,�ۊ+��v%��t;���_�ƕh��K��k%��~)��0��1��4��:���C���_��߅�����������c�x[?�å���ֵ��������������������������������������Ϋ��]\�   �   /    Ď<���3���9���6��5��1��0��-��+��*��)��*�݌*��r/���p��˭������������������x:�ڄ,��1��1��4���9���D���e������������d@���k��ʫ��������������������������������������ͭ��_]�   �   /    �j$7�;���<���:��4��0��.��*��)��)��'��)��w%��c��̮��������������������������t&�އ.���/��0��2��6��F���l��ߐ����Ǟ`���o��Ȫ��������������������������������������ͭ��a_�   �   /    �Y۠4���=���;��6��0��+��(��(��&��'��(��Z,������ۿ����������������������ӷ�Ǒa��r2��q4��q2��t4��z5���8�ŎJ�˝^�իr�өo�ή���г��������������������������������������ͯ��ca�   �   /        ��(l�7���<���7��1��,��)��&��&��'���'�lK/���u����������������������������������������������������������������������������������������������������������������������̯��ec�   �   /        �v$Ϙ1���<���9��2��-��*��&��%��%�،$�`<�qN.�wS3�yT4�yT4�yT4�yT4�yT4�yR4�rP4�pO4�pO4�pO4�pO4�qO4�qO5�qN4�rO3�sQ5�tS8��nP�ƨ���ֽ����������������������������������̱��ge�   �   /            �|)b�<���>��6��0��+��(��'��(��'�Ј#�υ$�ц&�҈'�ӈ(�ԇ)�Ո*�Ԇ*�Ն,�Ն+�Ն+�Ճ+�օ-�ن/�ۉ2�݌5��7��>��Z��k��i@���~��պ����������������������������������̱��ig�   �   /    ��C    ��*ϟ:���F���?��6��.��+��*��*��(��(��)��*��-��-��-��/��/��/��0��0��2��2��3��6��:���=���C���]���q��g@������׿����������������������������������̲��kh�   �   /    àNJЦ\T    Ô5	�G���K���B��7��0��*��)��)��(��(��)��*��+��,��,��-��-��-��.��.��.��1��3��6��:���>���R���c��c?�¨���������������������������������������̴��mk�   �   /    ťL3�i�Ұ\"    ̣?e��N���N���B��7��0��,��)�ٖ%�ϊ"�Ά#�͆"�·"�Ά"�υ$�΄$�Ѕ%�ي'��,��-��-��-��0��3��6���<���L���Y��dG�и���������������������������������������˵��ol�   �   /    ��F��{���k�ϭT    ʥB���R���O���B��7��1���(��j)��{D���T���W���W���W���X���Y���V���5��+��,��-��-��.��1��5��;���I��L��lU��Ů��������������������������������������˵��qm�   �   /    ��?��s�����d�    ��6شK���U���O���B��8��*�eI2�����������������������������͸���Q��+��+��+��,��-��0��5���;���F�Ϗ<��~i��л��������������������������������������˷��sp�   �   /        ˱d�������ܷc�    ͧD4��P���U���P���D��5�uN"��q\��í���������������������˴��̈*��+��*��*��,��-��1��5���<���E��x<����������������������������������������������˸��uq�   �   /        ��QK�א���������g�޹ZٹKI��P���W���P���B�ƌ'�\@+��s_�ǳ���ϼ��������������}@��)��)��*��*��,��-��0��6���?���A��uQ�м�������������������������������������������˹��ws�   �   /            ּq��������������h��Z޿NC��e���U���O���?���'�{S!�mM1�w]I��kT��kI��s1�ؔ%��(��(��)��*��+��-��2���:���@�ˋ;���}����������������������������������������������˺��yu�   �   /            ɯ\S����������������p��^��]!��w���Z���N���C��1�Ȏ&��~$���$�ϐ&��(��*��)��)��(��)��,��/��6���=��<��T�Ѿ�����������������������������������������������ʺ��{v�   �   /                ��o������������������z�޿Nt�����Ӄ���c���O���G���=��4��/��+��*��*��)��*��)��*��.��3���:��<�ÌC������������������������������������������������������ʻ��|x�   �   /                    �σ���������������������ג������ّ���g���W���I���?��5��/��+��*��+��*��-��.��3���8���<�͔?��������������̳������������������������������������������˼��~y�   �   /                        �܋�������������������������ܤ������f���Z���M���?���6��/��,��,��.��1���5���:��;�؜=��������������������Ҿ���������������������������������������˽��z�   �   /                            ��z����������������������������r���h���]���P���A���8���3��3���6���;���>��;�M�Ų�������������������١�ѱ���μ����������������������������������ʾ���{�   �   /                                ��m_�ܒ��������������������������|���k���a���S���H���B���C���F���F�ݩC�ǩ|�����������������������������ׯs��Ǵ����������������������������������ʾ���|�   �   /                                        иe|�҈��҈��҈������������|���g���Z���N���O���V�԰R���a�ʼ�������������������������������Ϯ�ׯm��°����������������������������������ʾ���}�   �   /                                            岊����������҈��҈��҈��҈��҈��҈��҈���^���S���[���p�����ɻ��������������������������ؼ��ͤb��ó���������������������������������������}�   w   #                                            紎������������������������������������������ޚ���X��\���v���������³���ʼ��������������T�k����������ji��ji��ji��ji��ji��ji��ji��ji��ji�   ;                                               귏��������������������������������������������������٢���]���]�״g���w�����������{�ܫO��D��������������rl���R��� ��� �� ��z ��p ��f�   ;                                                   ��������������������������������������������������������������ۅ���p���j���a���\���o��й��������������un��̙���R���D���6���-�ٌ9�   ;                                                       �������������������������������������������������������������������������������������������������������xo��֣���[���R���D�ۓI�   ;                                                           ���������������������������������������������������������������������������������������������������������{p������g���[�ݛ[�   ;                                                               �������������������������������������������������������������������������������������������������������}q������t�ޡj�   ;                                                                   �ĕ������������������������������������������������������������������������������������������������������s������{�   ;                                                                       �Ǘ�������������������������������������������������������������������������������������������������������t�й��   ;                                                                           �˙��ֱ��԰��Ѯ��ϭ��ͫ��˪��ȩ��Ũ��æ�����忤�㽢�ມ�޷��۵��ڳ��ױ��ծ��Ҭ��Ъ��Χ��˥��ɣ��Ơ��Ğ����u�                                       ������  ��      ��      ��      ��      �       �               �                                                                   �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       ��      ��      ��      ��     ��     ��     ��     ��     ��   ?  ��     ��  �             �%   ��  ��  '�  Y�  # �� �� S� �� �7 �I ?z �� O� �  B /_ �a 3� � � �� �� � � �� � � 7� 7� �L �l �� �� � � ��	 �	 [�	 �
 o8
 �U
 �Y
 �
 ��
 �) [Z �^ � � �� �� �� �2 �V 7X 7~ ø 7� [� � �) ? ?� �� � Ǿ � G� G� �� � 7( �, �\ �s �     �� �� G
 �(
 �         �  ��  �  �      4�      X�      |�      ��      ��      �      �      <�      d�      |�      ��      ����Ԩ  ��  ��      ����(�  ��  ��      ����H�  ��  ��      ����l�  ��  ��      ������  ��  ��      ������  ��  ��      ����ة  ��  ħ      �����  ħ  ̧      ����0�  ̧  ԧ      ����T�  ԧ  ܧ      ����p�  ܧ                      kernel32.dll      LoadLibraryA    GetProcAddress      VirtualAlloc    VirtualFree   user32.dll    GetKeyboardType   advapi32.dll      RegQueryValueExA  oleaut32.dll      SysFreeString     gdi32.dll     UnrealizeObject   ole32.dll     CreateStreamOnHGlobal     comctl32.dll      ImageList_SetIconSize     wininet.dll   InternetGetConnectedState     URLMON.DLL    URLDownloadToFileA    netapi32.dll      Netbios   winmm.dll     sndPlaySoundA  o~?��<�C��"C�ã�\<��;��j�~����H�`���,�D$0HUV�~-���W�x{�+��hT:<`J,ȸ��}D�3�3|$6�E4_tY	 /�l�d<�t	� s<�L�@�q3�u���c���}'>Q���7P�	�g9nLӆ��S��o#4���<�=S�1q,1�ȑsfDz��m���=D�rz����;�R���ދǿ£�+�.M�;h �@�\ؽ8��5*p0��U�7﫾��d�i��H-�����~϶�Q��@+�|���h94R�j!1۱���C���d���
�#9���M�8�sWk���҅�}�tj��S
���Flm��,��#�s���Z����R�V�9��<c���6�Ǒ��G����~�TtS�j�)��R$͉�"! |�����O�9g��%��o+i��'@}�iD"|���
:}�gUe�"�������ʫ��k�@��L�����j ��;�s|J!º�H�4�w
��%DT֡�1�P���̉(?�S���ꃝ�@I����D+��Y�qsQ��Ei��.2W��0��T��&;�|�g�s�	ԍULʘ�,�T�N��3$���s����!��<�G�
3��G�D�r�q	�dd9�+�·��:�9�D�����IP�����U������$nj��9�"{���$`w�
�b�%�ԹG�`�L6��\;�A%!�YU�0=�۫Ǥ��dZ��2RBu��ᯞ+���Ej]��:,�T�KD�*�+�2e,C�ɉ9 �
3�D�@#�L<��E�b��b�QcY.�yƋ�f0�9�Xj�R!g̉����G�bރ1�,�r�+��������7�����p0^�l-�N麺�u����J�+�냰0��o�%wI}��|�(D����
�����j{�r�-k6�C��Ƞ�@L�v������B���������f0�,}&��"�$�$��+"�$|��
�LD(�c�r"�I��B�9�$L���;�r����cuْ򂜈���k[�I,�p�t��_!W:�#�љ���F̙�@Y	
�\�d���뤇I�t�t�)�\W<L%Ϡۃ�ˍ��#�����,���|��N
u꾌;P�M���QTrz[_^���]��,�-��P�3PP!#)e�h��SV��W �F�*�	���W�jh&�6
������0�0��O�$���G����psRpj.��N�����AQPR�K0��V�� \���T��Of����S����7�P[�#�h��P�@T28N*+��� ��w�`��P�0pE4��J$h0�<�(;!���v�b��8�4M�* �b��;,��L	/b�@wЍ�C�{A @V8*d�����,��!�O2@SWVU�]��Lč�`C�F��,�
;y{�?V v�/b2�����&{H�$�sD����#ۃF�{����w��X/�oa2��P�Q�F�ߐ`�N,�1�+Kj@3 $Q�7!�0�'V����r�����d�(@YU$3����4�������QFGA�nt{����͍��DuR�: �-���W�t�R��h2Q��11P?
�L&�A�R�?�aS@�j�����H1�*(7H�%�uC�K@����/�P+4��%¤��(�W�7�q���"g�;h�F�]^_[�Ui������@[���?�HXX	Q����E��\V�(~�r�X��vtR�~�ÿ2u�D3"�Z���X�Ta�uŚ�����Т͉�f�MG���H�~¸�)������V��x\��>��`X<tX
��0P�'. �U��FX�Ƈu}yʹL����z{l1M�@^�6u�;�}4��F��U�,���t��Ȋ�u*;:�f�����M�����0A��^IY�Ft5;u*X0�����/x��QP�9��4��f�vRP�3��0Y�I	?W����V#A���'�Pޡ�CE툲tdM�s�^}(KN��!��`-�}��({g��R�����C�Zf�`;2�=2���
u���B���G	�QRV����֊���1�}�q&�nH<+�)6�Q^2 ��|`ʌ��H��R�K�K�3�/�Q~��`��@qt���F�)A�6��n���Zk��;}�u�(���'@���XT�ss�}+ԜI�^��N�E�@�-�-@����,�Q�]4�9�\���t$n}CQN���~���!{@PWQS�ORe	H��	���9s�msvbˬ���AE��-�l���8�F����bNA@��b�~�Y����0N6�N�cH��Aɔ�}�U�ҧ��f�*��n����
�tDRD��%	%�#j���XM�.A֞f|Q@e�IZLhl5oM��$�Td��Q����ʄ"��o���*0+6����;M@fA�W�6�	k�:mYP �EA�@<H �|��'��,��`��Q�vP���`:���P��t,x�QY�9c��e��+)fz�"�2�%3)���ϚJr{����h�-���V4�o�LH��Ap�licaton erǷ>�} �u��.�The��;<c?d��%s5�l��n�t�b��a6nid�SDL�G53�d,al �+3�*	W%'c�d�us�32MoOagaBoxA�wxtffk8��l�?ExitPI��L6C�hHand�Op�V?G�tM��Sl`|Virt�F�A��c�M��vL��	�������m9ӑ	�"PD<H�0MzI1�	���]�  `�t$$�|$(���3ۤ��m   s�3��d   s3��[   s#�A��O   �s�u?����M   +�u�B   �(���tM���H����,   = }  s
��s��wAA��ųV��+��^��u�F��3�A�����������r��+|$(�|$a�  ��  d  h
  (�  ��  ��    @ ��  ��  �}�`���� �A�T$�R���+ʉJ�3�øxV4d�    ��USQWVR��W �SR��j@h   �sj �Kʋ��Z��PR�3�C �K �C�K�KʍCPWV��ZXC��R���F���+��V�K�N�׉�? ���KZ��h �  j W���Z^_Y[]��    �`  �` ط` ܷ`                                                 `��   � �    ^+�Xt� �Q  ���s� ��3�D�g�   �0FZ���	I�g�� ����|9��{E=ܠ�򹿂�����ıq�~w'�j��5�]�|&j@�mz!�9�������N�Eh�r.���5:��t�_����v� +��4/H������3��,��Fw�ʏ����8��Z4�>%%"���^��A�I�[E��B��VAy�Z���PL��Ѝ��`R��#�)�{� p�n��|��F�w��sx����.�Dq|�u��lm�R�V��vm�W�m�:�Js��B�D�m2´)(��Y�O0�鵅�2�8m3aV��z#ٷ�f�1�F�I}��9?Gȷ�E��v��~��,���ڜ]k�ڹM��
�� �C��������%G���?j�9�=R�X^Uի��D�1YL�qP/Ƭ�?I�KŸ#^y�k�M��O�F�
�j:r��g'��t���z�Lt��t'a�a�rcY���h�vM�/��`,������'�nq���m��8��&k�ǉ��!8�XޕE��yr���;�LE�e��OD+���Wڽ��]�\� P���DT7�a��͖,`���_�9
��͈�t���I�%�B%x�{�7=}�;8!$#~�Co�����k�d
�AB.��X�0w�=���v�#�-� ��)��,\�&����ZUd���*ct�I2�[C�M���B�FN�	���BC�Q�qJ�K�{�d�"��ٳrQw4��aJE�^���e�u�w5N��bk��J=H�fx�����gW͙n�!<C�O`��eȁSF�x��Q� \A���L2I�.��.��"�� �h�#/բ�����1�U4)��*d?��5�UL��̙Z��=X���a���)_�|�����P���8Ӿ���xS�
�v���`� =�ݒ�$�����,�G6n���ƍ�Q9T�iZ�1���M��N��H�e�
�%{R���`��le*g�t���r#|1����r�o���oV}�s��ꁈp��x�R�������oa<�����_g�r�o���=0cqb�=]�W�Y�_�]�K�>�@�>�4�J�H�2�L�9�+�1�+�-�?�9�'�"�,��$���(deavT��(���:Ј�'���b��1�jT��A�u��u�+�&*t�6�b���҃("Ny4�ѝD����^�F\�m�O451l<���I֯ c]SD���D�)�I�D�>�p�D��(BO^KWG0Ѥ!����?�[V�R3�`�����;�0a�����DW��7�e	��0���?���є��#���\b�x�\5����Y��r�.L��n7�B��ׇ��^����GO��?ic��m��>s'��Y�hp|�֢���H�y-�G���
}�ۅ�<�:�[F2?�q*U�I����i��O��w���փ���0o�<����G�R���=�Wnh�\ϡg��C��)���,���%V��|���:���Q%3;�E�_�_�@t��-]����|���j�h��;f��aٝݏ֐��b�ܡ��z��D��([������������X#�����R��B�l�_��%���� ����MpLF���e��Zm[��i�#&���ؖ ӎ<d� ��qԌ�o^sѲ���� "J�b|	��Y�'��`��l��o8��Nn���g� �O�+̦-`�6򒼐x,W�ܢK�UzALW@�
u��!����zqB��n}_�� �{i��v�Жd��@�96�h��ɳRܻ���*���V��+gq��T�w��13|�ñ���i���`�����,S>Z����_���*Q�׀-��*d5�ZP�3�}�᥽�N����k�N$���@��w�f,��H�n�wMp����x��6f����,�C6��!���i�Fn��ʯ�K�����b�P��
����,�O�,��[W�6u �%^4����(�'7�8A;B���4�����L���.��'ek�-�C*�������r��.�g�FY������i��'f���#~K��q/�)�eȮd������$xŒ��Ԟ�̩W�;}�w,|��t0V# j��)�����������m��4�n��|i�F��NK-�F�)� n�����IRPZ)1Ή��_\sp/����WW�q��jOlx⦨�Ԡv�|P7k����m�6��~Q�?�g�7Sm�&|��Z[������P0�Y�]���#�Fo�5%���E�N�h;���C5�/rjc����H�`�{c83���EVf6�߭:�ga�X|Ψ���TD��L_ݒym�ә����Y��b.�1D{�,|��k��%{-e`���v�kGH�,t,	C#�2�l[E��@�֖�H?���޽��SL/e�$�=���t���sߓ͵�G�0��G�fo��[I��/�&�(��cW����[ �m�ڟ�x�9��E�g��O
5����$�p��v��X�]f3DNBL�T�Ɔ߂�#�jA�T�����i���S�>������9u �J�D{vXW��}LWZB3�0�.:4^���4P!�t���8��B.���4�B����$����w&�7������wO�G����W��B�vu� �,�
���5q�J>kC�i�+�:���ߟW1�����uo�;߽Eּ͑ta�-�Q跉<��*ӥ�L�Q�xX���g={<��Kz���6����vҢm(ъ���Y�(c�Dz���6��.�A���w�WE\�[D��pzo8A *�N�Aʙ)Kj"�sS5�'Eŗ����E2�{\�[���\UU�J*�O�{&�t�:�.�OBUJ���|e�:���O��v���BH���/B��P�`����R���)y�!��Wf�3gF�PJ�_$b���,=���)�$��W8�t�p�12"5o�<P�x�'{�O4~����aBm%c��vƣv[��/��u���Yg&L��_�?5�H߱.�	�n��Qg����T����bUn%�cVZ��f�-y���/W�_}�Kt��5�i�>(G�m�\���r�i&�?2�c�x�&��z�>�dt8��:��JU�6���(�_,�3^n�:v�&�({��wWR�se�9���[�ư4�B(q���y5����xdZ�nO�L% ���y���������P�(�8yx|�"� /~\|D�;E���m����nK0[�j�P���Ҧg�3\>"��\:e��Ҩ���{\�`H�.��s�N�q[�P�n��զg m�8��s vV+}����?H��b*͏V���t
��aX(�/P���tCv�&Ɉb��BH >�����?�_�9M��3��B�pUx$�,)9��D�{�$Ԋsa?��N-�La���9����3n���:S�[u��`��q(��E�̝�E�Ӱ�\?���FĈ�  �s�fÆ���SŴ@Q3�(���2�}+��ؽ3o��7�U����� w�'I����_��1�[(�����x�N�N�:�&����X��_�g��y{�!㋭7�W��D(�ZcŘ8:ϼ���U�h�M�i�*/q5:{����bP�qi�ްGP9o����%�*�z'W���'�G�|��C��6�[u.�=�>ZvΨ�v�@@	��b芻v%���{��hp{䴺�AK�d�COe����E�JԎ� �Z!�m�Ԧ7�'M���Tm�5�h�VW�~�VM#�Rs��Wlę��QJo%��b��'�R����㐀�u��Q��c�TF�w<˗����Tz�U�Kم��	�b2Ό�,�"�t~��Ki����j�z�>�Dh�Bi`e��
Gp:�-QOʷ��ei������E�CT��G��҄J�U�����7�[]DUS����C8��S�`�����(�aA�����������|�Z����?��HQ"�#-��ܔ������a���&����M��?&0�|��=AGv����T���*�J��N#��B�[=��Z�� ������Vs{�3�/ױD�&4�JD�J5�,L`����Hdߜ/��봊ǠBC|��v�_�S_�4J�bT�If�vp��q��rq�>H��v��I/`,TK^���Cn��z��ܪBW�t�0��N��>��0.Ԟ�,�/�����Y1�}r�*�ZKW��/5��F~<��N���_q�c��8p��]�Yk�q��eD9V���}��+Ӭ%�s�`.�R���b�1)��tK[ h碻կ��4�0�3��'�jԏ��v��y�`�/����ڞA)�bE�`ʅ]�����-�����ͺN#����2�L�n�u}��� �+t�R%H��Tċ�`�ů>P�#�R�"�����|-��.���Vr��n5��B�����q�l1��I9|�w�&�⏜k�����M���a�^��R�I�l"H|.Z��|�9b m}�S�KKN�ծ�N~�-����z�W��vB���n���B�#�d�+4l����j� O,wԍE$���Aٕ��Tk']Y4�C탻����o���E7Ҵ����ȓ Z���D#�S�e�	J;�I@��,b��&�RO�3q���}��
��ῐl)��/�kU��L��� Д�;-b��@�~<	矤��m��J)V�.�i�ĵ�G&.HN��W�w/�ڍ��C?}�%�^���=���W��-��9{"��^�Ԯ���;7��)������>�����rZ|b�e)�Xx�}F�Kx�wJ"���8��=:�W<ѧǸ�M-yx�G���g�?�Ql���Ğo��\C�d�C�X���m��� %F��0�;��S����uк����}�s�|�0z���<��Z͗Yn� Rs�㒲�������LEBIԭ�墒�#�����W쑒Z���\;B:&^ .{�pZ@�o�V��ak�A�VO$A���AQ;6�6Vį�UD�79л��0�+Dk�ŧqL��*�#�c1�zy~��QP'K���E���2�z���Wy��W����a#KpEm�aQ(ܕ��r����ݲ��^��6j��n۴V�9ޒ]C%6�N�1}K�Ӥ79�1����ʴ�K6���~�h	�`$�I�k��w��"�G%�� �"w��IN[Y��ͭ�8�6¾��Q��7k�����z�z�aB �,c1[���.vh6꟡L��P���F�<��g���O�E��	ݳma���5ۜMJ�o��l/E�ˮ�P�Z�Ű:�� ��.���;4�${\U��I:	+�Hn����_i� hm����N�R�$�3=�T��à*$C3���h� ���ʴ-p��^�[iÃ�c�;0�2bP�v]�BzD�J�RDO���L%�_؟aObAj:C��M�ìw�����.��G��ޛ���q�����v�j"���gWG�ҙ�E�'JN>V!^��YMh�������,a;e��Jz��@�s���A_��{fB?�ъ%��;kv}�h��k}Dڥ��%�Md���,�)��.C%��� (?s_���܁4�0p�|�c�bi�Bl��/��^g�Ye5���Ad�y�C�U����Qc�n�v�2�zm^]��FK�+ap��AMz�%x|�L�z��7ӃM-�7#\�W���j�f���"�,[�!��C�V��a������<��}��k�W+���� ���EG�4��N7yK�%~��
I�?]�}>2k�o<+�Ti/����K��I�B큵C���bP[	b�%NN�e#�|�D&F���6r�pޟf*,7D���BU��Q�Q������S���.*��|�qݤ���#�������@�a��9!��yk��1܈ۅ�O���1�g]��V�Zo��)G{��W4d��$����{>���d]�X<+_�E�)��o6\#������v���N�U�Rj�Ш�TZrQs���b�#��? &B���p�7#�^�� T�s��N~ۦq�h���� F�iU�����m�'L���ög��5��[�Si��Pw�ZD9��F�_t���?������fk�|A¶A���N����\��OQ���`d9�Ψ��%�5ȅ��k�����lAv���D�oez�|^��k�-(z3��e�'��Ћ+��(3�
�Nb�S�L�G�f�{9.�Y��5E�EY�a����Ө��*ܥ�O8/��/Zt���@�$��y*��Ő����)��7�*�=��4����K	0]?��}�Is�h��
���=� �Cr�W���C8�𚭉�j�����3)Z:�%ӧ���8���/��RF��2&�G���������H/� ZH���B��?|�s=/�!L�ws�U��{p���I�(�T��1I�9N)~�YZm]���CH�Y�\%���!��~)Fp��� T�K�r������m�Ͽ���+ ��e$_w=Hʺ�l�.T�s���n�   ���   �������;   ՝cTfG��\x�~5f��C���H8g�<�Ժ>rV.�bߙ�C�i��<��h�Iph�r�	   ��   �r���tØ3Ð`�   �d$�+�d�2d�"�����u�#���   5C�^�   ��sR�3��r�+�d�^�s!��`�   �d$�dg�6  dg�&  ��$   ��s�� dg�  Xa�s��s�    �� 3ċ$X��A �u����8�   ���   ��Đ����5h1p��_���c���r� �����U�5S�ȁ�H�5S��3�Hh���W^�� ���k�!17�����C�   ��s!��p�@��F�J�����u���    H�y������a�r�ê�ݴ[�g	 �G�O��]#����3���+GJu��z�Մ��C$�و�_�8ʪ��GJ��j�RL�Rks�����[8��A���?�l�H��
�:�'��y�ǲ��T7�w��]@h���    �,$7  �d$� �%���   �SA)�          >�  .�  &�          K�  6�                      V�      i�      V�      i�      kernel32.dll user32.dll   GetModuleHandleA   MessageBoxA                 ��  ��  ��  <�  W�  |�  ��  �          �       p   �        @                 ~�\N^��2�J�x�Ws;nn����g�)�'/��W��o�
lY �f
��d8��RW��hB�H6�� �w��e��l���D��H-�^]Z�]���b?-��I|�D4}���h�����K|���}:�I P���?�_�c�1���v�yw#�O����w��r�Q�1ա�G���Uo[����            ��	H                    �!�=�P�F�>~� %M�:v��ō;x��ӨS�R�P�(�{L�l"K~D)�HV����nx����s� �7�'�>Z�s"i~Qm�Oώ��qZ���� �%�$�f�}J�e"thV9�WV����{\����!�=�p�.�r[^�occxK*�[V����~
����$�;�5�*�}_
�ne'p	�vV����hR����6�=� �#�mW� gucJ?�:5����nI����:�7�3�(�{P
�hct1G(�TV����zR����5�+�%�4�p�s{te@ �0����{^
�Ȱ�6� �1�*�|L�krhxK9�����y
����=�r�8�5�nL�rcj0%�N����e����s�3�<�"�>j�s"AxI(�R����yUX����5�7�~�L�{_�n"jxB%�����lT����6�$�"�5�wP�cvn~Kl��^f ^6QJĉ	�ԇ�  		
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         